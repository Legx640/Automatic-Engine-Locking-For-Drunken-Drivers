PK   ���Xw�x5   r�    cirkitFile.json�]m��6��+��`��oz�oIn�p�\{f�^w��ؽnw&�`�����EҦ\��� H2��Q�X�*���g��f��6�f�K�}Znֳ��OŶ�R���g���b�Y�}[<~�=�n��~{l�r�u��}/�D�U���d��Q'*je���P2��E��g�?�oG`d�x����9P� s�"�I�@E��́�/2*B�H���"#s�"ċ�́��m�P�!4����JF7�d͂n.���`�!4��$Cht�I��,�f��Y�'B���N2���趓�Y�m'B� 8�t��鶓�Y�m'B���N2�fA��d͂n;���v�!4�� 7_�m�-����|�Y���7��Iý�U�Ϗ�u��-��iX��(Mx��X�*�ZĊI��*:N�1Y7'>�׳�YN�('�|�38�ء���%�Z�D֪�RIY�Q�p�eS��d��S�zr��9V�Pv�.^��VvPv�.^H��$VvPv�.^(��VvPv�.^$X�%X�A�1,�x�be�beeǰ��E��]���ò�9Vv9VvPv��$��~58���c`~��X~���@���`��#,?�g>׀��2�������8���c`~�X~�hˏ����{`��#,?�g>K���:������
�8���c`~�S0X~��ˏ������38���c`~��;X~��ˏ����`���p�?q���?88���c~�Os,��nˈUɒ�Q)�**�L�2I]�u�DQ�C]�����K�U�2��*���`�F,e�FiW	�Y)EmV�ee�7��
䵁#&��ͯMREe3�k�䵁5,?�
'{���1��h8<∡������C,?��w���+o��%G�X~�
�ѫ�N�y} ��pm��es������S�\��Ҵ�#�Y�<a��E�D]�i],2ϝ�:����A݇��Gv���}�{d��
�݇K�Gv�Y�4�����q��c5���D������OTZk����D���;��OT\���0�����Ƣ���)��1�ތtoF�wL�7��[�n훖�nMҴn���w��t��V����D�bm���gl��&�s���m�a�!Fx*�D�N��PÄaʁ@�'p�E
���`R�����pk��
��OA���)���:�����f�P��ro���}FʽI#��R�ix�N`6�)���!�'p��
�1�
�s�B���J��Ha���Cn��Ri��"�4���Q�m�$M\dL�:Vo(�Q���"Ds����az���e�u�EY�U���L��"����$K4**Ĩ=�o>��%H�|�6P�	w��N�#��w_�[�"��f��ҋξ��?���@ԙD#Pg)1�@@��0u���X#PW��ԕ)�0uE1�@@]	C#P_�d"qVg�av��7
�/}���f�QH}YD'��f0�B�K&�8�l8�qR_N�	f�9̎���R� N8����8��qR_��	f�9̎����� N0;�av��sq��q��>$�BN���P�n�*��]����ʲ���$M�m}��5�܇��\�����a�:���\�"�	��Q�r���]�#��?8*P�Sp��7b$0܄G�u
�vaG�����@�N��.����p(�)��!1�o���:W�X$F��kpT�\��j�y�S1��� ~��k��Z�xX�l'
��`�C��E�v��k���xX�l�	�&a�_��E�v�l��ږxX�l�	�&a�{��E�v�Pl����xX�l�	�&a먗��E�v��l��Z�xX�l�	�&a먳��E~Y�&.����')�i�I�:�s�a�����4q�U���4q��-�;�4q�U$�i�2[�l�H���*T	�4q��-D�v���4q��-io�H"�i�2[4,Ro��ˬz� !L�9�Bd;M\f|	a��,���*�.0��$�wk��"��o�&��ƍZ�����}�xV���	@��_��Y]=�B$ %�h�g���0��m��� $���]c7T�D�`t��Nն��9f�Ū9��uZ��8�����22[�����)�V�~(V�UI�鵸�U�(0{-N�RQ`0Z�ۙrCuB��-Wmqh���Vh���>ch�@ ���)�j���f"Bk���ձZI�ru$�ջlȃK�]�V���]���]�r�k��d��\��� (��X�����ve�,�6�&)2�TqM����f�T<�򖀢��]h�1#ݢ���ba��(����wZ���D/��vŮ�Z7ϻm�:�w[A. P?6 �@@�8�0�c�ԏ#PoK �@@}A.#P_����0�� �@@��\���8���f�QH��\N0��`���/ȅ���f�QH��\N0�`F��/ȅ���f�QH��\N8����8��qҾ �̎s�G!�ra8��8��qҾ �̎s��!
r�Q��9 TGA.4*��� (�)�:
rA$`��G��:WGA.����hT�\���(������
��\� �V�Q�r���� D�
~4*P�Spu�H�Z��F�u
���\	X+�Ѩ@�N��Q�"k�>(�)�:
ra<�i.��Ƈ�&䚄�� )ۉ®i�.��)�iB�Iغ
r�a���&����� )�iB�Iغ
r�a���&���� )�iB�Iغ
r�a���&���� )�iB�Iغ
r�a���&,���� �ea��l���\pX�l���&a�*��E�v�Ob��ev�+8,R���e��u��"e;M\6	[WA.8,R���e��u��"e;M\6	[WA.8,R���e��u��"e;M\6	[WA.8,R���eAlo(�EG�御 ų^���\t��r	.�EG��ų����\t���
r�Q<+�o(��:��b�׷9\ ��v��R� ��a�v�[
r�F�}��n)���h�o�-� 0-��L��  �����䢣`�\P���(W�SpA.:���\���ru(�hHy1�{ݫ	/���(�u�&� ���Z�����r݅-�EG��@�予\���r�䢣�r�:�������f�Xֿ���Ͼ,����qUTM�X��m�lg��S"$���8w�;0�D�l>��1!��2��U $f%mGy[|��5:YGI�x�8���/ʭ����?t�C3�.��@Hb�~d#Q�nD�B4��nD[:|2��%��B�h���toRu`N�7'�f�{{�yhd��0��x�yM�Rr'1������$���on�G̤�4�ւ(��up����R��;{T!03@��.f��^}$m��xH^l�ϛ_�zQ�kW"�f��ٌ���oy�����O
o�Wq�c�W�/�Mĵ��|pi����+=8=E'D�R]$�*�*:p��"��I]�)�3X !�Y FhψN	6A,��-��61�+����� ��8:rV@���C�h4����M����c'�WI\����Ȅ��$���|eB��8
��f�3@g[��I׋�^#�J'@L���	1K�|ᡢ�z�Ya�^#8{���_��y�>�y�����i��|^ր�3�|o;7��/^%� C�_�,���Y"2D���Ȃ�/�%� C��^Y�!��.�,���Dd��DK"2��K��BXO���O0�t��	�T � F���?���`G���1�'NRy l)S:��dI*�=� {J�؟ I��G)��r�=�c�O��� �S��t��)�T {�����?��`O9����%3�x�ߗz"�u���������*K|[VeX��c�9Nr������*K||,?������� ���s�H|^��+"?,?ǁ������ ���s�H|^�F+"?,?������� ���s�H|^��*"?,?ǁ������ ���s�Hu���0D��P�]G12�G%X��#���C0C�Q�@@�������B  F����u4!#CtXf�:���!:43t5������bd�Q�]G12D�)`��#���L5:N3t�������bd�d��S��������hJ� :l�OǣJ ���E�I��\�^Y���H�� o
��m��`$�y�]��DJ�3��&t.�ȉ@D��xT	�"��@�	Q���>�*t|t����J������Ў��ty���K�g[~��}��>����Z<����wdk%����
ڑ����#�[+VG�݂���`t�:������ޟ�� T���Ɍ�j��1e|M"˿��>ko�G*
aO2�2n��<J5=�u<e�����S<i�#=���%<������ ���bA���->�o�$��|� .%�9���Y�>�o G��e�/�=	>���FW��}���V�!}��C*��?(պ��ܾ�2������c���f뷯�Y��~z��|�� �7[���3���^�o�=�o �1����<f>���f�<�У �<�4�L�;ϸ
>0�a�O	{���Z�u>{�Y֦"��2%�B*���3#1�fě�Ef!��q>3cܘ!3�Ι7k��u��rg�鸛����h�
�����ɾ�C]�AnzpӃ����7=��!�y�����ob�^ng�0P��4@�.��1D�N:h�z�Ui��&-�Es��Ӆ���sh'�����C;�D G=ўJ�d^�|D�O �A�h�_nrosr����3��]7�W:,�v�)t�����
��H=;��!��g��:���Da��Ϡ��&YQ���SBY�O���6��^��:;L#���gg�iv�#�����UN���2�Axv KxoԳ��$�E��g�(��K�k~�-VE٬L46���2����-\a�K̾����}I�/	���_���d)�/��K�u��3�=;���}f�g��� ��Zfw;<��ˏvה���v��L�-v
sH���9hn����4�-M~�&w(�����G=�&�T�V��BZ�u�Y��O;3n�ƈ0U��g�����:�U���:��)�X5�ΌԷ��q�>�G�39�߻��m7��v�lL�M�E[��n�Y�:&���,穚G�n�^������И��Xk���.�F�HU��Dœ�l[�$�<��Ӵ1�}��f��݄�g��ӮXW=PP�o>�l���Ξ�r[�����Ob~oX�\}��OXz���D�[��^���dJ�y���4}Ҍ'���M�����{����3�ؽ�7:��������HJ�|�m�kcL��g�wsu>��X=��}k䚘��^j����{������{�;{h��S�/>5ۿ-���9��m����6Z�;��=~.��mQힷ�lR?��f'L��� &�*�w*��G��$c�\��v�W\ԥ��V���T��Q�zz�J�IU*e�^假z�]����R-�gÎ�g������l�ɠf�9Z�i���D���4�����-�4K�n���}|����Pg͸�����*�2���8I��I���p�&2�5~�_����z��kif��x-��Of�kB�1��~.�8^Kmu=^s���CG�ׄ�*����~8\��{7���z*���fU7���:K�a��a��fW}�0��-��2nkV�<ESFRf2�Uɴ�Y�ʴ�Y׾��q��&�?w�W?�}��+^uT�iI�DE���j�WIR�q��5�?�'�\���QZ�I$���򢬣X�YYdE����������s7ͷy5�U��I��yUFU[�MQ��I��O?���1�2�p�^���O�U}���E�eEi`M����<�j^��YT���L���f��c�>A��jY*���Z(	�IfHf��]�;P�_m��36�A�\��U2��y1i��2^�M������s����b]7�����o��U�3��,���Ǉ����z�u>m�׃��^y���m�����u������U�P���z�`�֯%�,J�l5�RE��1������y�7>k�4ce��7��%�LEy�ga�+�=�8/c��Um�U2�bZ�2kY��e�P��m�4�^kU\�Z3,S�eR�g�$2*�XO�mQ2�.+X�����Ͳ�{jvϏ���w������ӟ����~�<o�+w��ݧf���v�����n�]��Z���O��l�8�����m�b�ԫ�N�z�?7���u*ӱ�:���z�����]t�2=s���
N�����Һh����ݏ����i��j���$�����A��d�:uJkYs%t�R�ڡ��8�*!ˈ���Z���u�4�s{@��eݔ�bi�܄>���a���ܢ&���:��Os��Y��oʥ��r�i��0��H�`L[�5�UD�Md�T��sTR�z�h��s�C����)��5c��õÝ�D��I�#�jpϸ�)��I�Pt�?�7��i�
�;��n�Ș�@��ӣ[Y�N�=�T�}T$t;�uk{��45`�7���]N�_�6pŴ=&�}�{.�TB�Z_j,n���"��4�YSDU���������1����@d�1���^ƙ�������࿈�0�[�+��l����k���vhOγ&�D��ɢ�e<jӘEeQ�~�ڛ˂�'h��P{�͗��?,�u$Oci��d�r�����ZH~�7����y$�r%ɏ��+��� ��/W�ӻ���o����'�i���V��]%��'3W�/���k+&��H�D����ʔ~[G��2jҺl�v	��t���"JS��3퓥�hR�VA�&h}a���ݥ���V��!�Χ�O��l�ެ��uȹJsѧ���5�26��S��F�=�\;"���btfJ��Z�ʤѿ,��'�feq|�dړ�?~j����M{�:��� �,�-�OM����ƻm�����e����~2�8~7�4� �~0��E�lw��}x���>�]�(��z[|�IU��y:����z���}�u��af>6�Ծ3~��������w���h^�W��$�i2w�˜�cW�}��a�U�ҹV�,��;��
Ԋ�X�Vp�V8َՊ�'2vE+�virϕ�ݹ���i�fv;���MgM���-I��gcWF���j^����H=:�x��T�V#=���̫E/�qG���ܭFq#��!Ո� =
[�֣=� EAo�"��`NU�m�,�ڎ���0Ώ�털Om�{�ԩ���Siض�T�n�JGPN��#5�KԞ)��"�v:8p+.��]�9J�v�@�g��$\�Fp*���XۗU���	����^Vh�@ㅭ'��x��>`bXr��B/���*4l���s�ڝ�d`;�������ms�������[`G�{�c�Q=�$��w緵˙[5�$�-��V�V�Peʁ���ʔc��c�)��J2$��yN����]�2�Ӣ�F��ܨћ&�!���6~deJ<g�$��<����tK;ߤy��j\�@�l�\��,�䠍�B�V�+�m���)-Xh;�`"��]��ɔ�w<�I�u�J��&zdU��+����v���O=\ʪ�w����+YV��q#O���a;_<8�^���+��m�?�:�J�u8�0��Z7P|�'��v��i���vogݰ߸�&�����Ew�uS���A;{R�v��(�ӺT��(�
H�1
,
2��s0Fc�T�����v\����|`�B۩̭"��N��ʄ�f�Zq���iet�*���^y��{�X���#�Nx|5Tɰv�|�	����̣n��3�+�3��.YՎ{C�ek؎�ס���$EƓ
�ia)���K`�
�0�`7V�^�7��z��&u�>9K��d	��)
lw�C��;S��v�ig]$�2s�ӆ�˱G5<[�}�'+��djX,�n��󏠆�͛����S�^,h��LGB��U�l������T��[�.��A�����އ�#��qG��<�����ӻ�:7���q汇ƾ�ɕ%{����4�;�G=�#�ڽ��d
�*�Nr0p��wl��d?[|)�a���M���I`;�ڟk;K^+�Ɛ�UM�j����w��%�r�sg;)��dz[;_k6�-W��ڿ�f�,V��S�WO�_����)������w�gS���ǯ���PK   ���X��(��8  �8  /   images/02932828-f6d4-4923-89fb-67d65ebd103a.png�8!ǉPNG

   IHDR   d   �   ���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  8kIDATx���T����������tX�,�(HS�(c��5�ؒ�1&�3��&�F�1�?1Ѩ�1��i"(�.,�l�;���o�웶�]��|ٙw�}�s���<ߘ1cZ����&�x<��z���K\\�466JKK��=!!a��f���f�w||��{���!x�#��1��|>�< �\�r���>�v�q���͛eӦM2e����dܸq2l�0ٹs�����	��}�G�ĉ���J^y�)//��=�IIIr��'˜9s$%%E;�0ٺu��q��.�E�u�(<�]p�:,��g��:9##C$999�x�m۶Iqq���Yd��=z�̜9S���Z�߿����K����g��C9������'//���'�0s:T�-[�_�y��Jee�A<�~��f��ٳG.��2Y�~�����KlϧO�>2`� IKK3g�޽��555!�A��Ғ��w�O��Ө(P�6rݺu�t�Ґ���v��an�U�J�ٳ�lٲEv��%EEEf�u���Y����3�\\��� ���s�]�}�v�����3c�p�n�4i�2��Z���^�>r���J��/6���gAX��t�0ax�R�%J9�t�$(u���Pޚ�������_���:�\��B���w������a�\���ZxFvʆ��n6���q};Vw�%��W�^�JAAAȯ���S|���c�����#	z��!cǎ���z����iJ�=�!v�#F�xAW��M�� 7ʶ}�����o�'�|R=�P����
�%tvn1+Y������� �畕+W�"L�n�,�e���V�Q�������ؕ�;,11�E�[��r��p)�*�B	��-�N�����P�W���9~�m��N�ͼ�_�כ<���
-���?�8O���h��TU�.��w�q�lۺM�9��y�	RUY%wnO�
As��>عc��=�9����o��V`��+������J�,^ I	>y��G���e��r�7N�Q#�ˋ�?+�e%���$��		�fa(^���_���%�w����7r�5ט�7��>K�K6� H�6;D���}W^ye��gϖ;���S]q��΀Ҭʐ��������<�w���eM��*�q���Q�Ƀ�Յ���&3$>c��dű�;�H�lʢ��d᧋͹��\I���y���/iƙ��v�_�w�<5w����J��������7�IrS��Iz��́����n��{ｆ((ʶv*�W�=�c��y<�ET�3�^8X�A�W�ҴZ���:�h��47���5�����|��/���S��رn�(���o-N�#�:TD{P$��߷�rK���.�j�>S[[kvKT>j�js�bn��|<����5��Zb�(��s�D��Ǽb�]�yc�ӑyU����<+,�9cΫ�dT��?Z]ǹ�����;�4�n��V��+**233�#��i���|�8��$:�#���A %H��<T� ���Ȋ��KmE������"i�x%��@��;\�S�Ϯ�x�i�\�y� q���)��=���|�^�'i=�IF�A�OT6�����2���U��%ez��U��KL���C$C?]��MQ�G�EM��Ç������޽{�sss�a���)!��Y�Ǒ����=?p��G�e���u�1%T��Q5���]��SZ�S|2�~)���J�����LK���ee]��|��t7T
 �-�d�s7If�Qr�ٿG���mPB�{�ϲo���'�Jz��뽪*��I*<$���Ȁ����؅�����d�+wI��)2�?��l�����3Y������Œ���z�U5��a^�T��e��ߓ���"m[D��[�r�jY�R�}II�T�6��a]��t���O>	�!2����������<�4��q*�.S{dȼy��;J�/QJ������L헱��K��s�qSJFZ���`�������u�����oB�C]���RQ�.�L+�Aj���ŏ^#Ǐ��+�"#�$9)^�A�U�2��5r�_~*{t�#ξI�g�aW�W�H�����#��Z��m�+����3��"��d�jƏ�"%����ܵr��W�ލɘS�	��V����by���� /��1N�����0���s�ƍ1-��7L�q�5*;??�:%�uF�c�~���F�t�l�ʽ[d�?����)�~�̙�A��_��dמ*��'��8Z�N*W^��,zl�L��{%�N7kX�]@�ؚ�BY��������՗�nvqCc�46���3H#?�l�����e��"�}kP��Ƹ�V�;NO�d�+��;gȌ�#���IWs�ޯ�k�3S���'ɱS�ɅW>*k�H�Cg^e�+7��P9�}5V�}�,|d><�-�!!  
��+d͚5F�[�X�s�GV�p�\|Z/��w�HUu��`���x|�Kj�z��F����˟�8KN��aټ�e_g-��Y�>W�x��?#U���t����X��#�u�����o�>C�\����͑�+���#�}N�+e�[䞟-'��_��o��]R]� �����>SN��)5Mr�n�� W�����Ø
(F(EVku+FQ%2�V�u�r���l�XR*��U��g���푕,�Jk�fq��J�F��x����صߛ"���w�a���(ݱN�K>Tb|��Pb����݉�e��WL��zD���}^e�;�͑��r��ce��RIJ�Ib�W���o���
��/c
�ȅ����T&_pgTcֺoX�����m�H�ٴy�"����2u\OeK�RS�h��#E�o.uv���2E\��x�����c&��?,������
"�UVP��C9�l雗��v�Ab,ئ�n0��:i�yґ����[~��RY�M���z�{?}O������ҝ�7r#A�aR������Fe��N%��H��
�%�>?�(�����!��&+9';IW\�Aۿx_���K���{fF���U[H���2�G��f)��kŋA~Y�Ab4b;i�A ��/WeZ�N�8:b��F���)���Fz�<��&��Z�+��jw��8�i^��=UR_]*��i��ϙ ����M ��� i�	RV^�ȑ}5F{q�0��y؆�����o�x���vC�r�Ttb����j�So�[O�Yţ�L"R�qd�e���wX��7G�����;�c�9
�)��l�X��I��'����d�`w�d%Ii�#GXٰ��D'�V]S/{�5J^f�!�X���Ȗ�k���#���Ęf���� nϾ��̍�@�y�{J�^�r��CU��5;ο�@�����/��+�T�iI�Ĕ���q�All!�66�	՞�gw�1I>x�ߊ�:=��	#G6nq��p��~=�)�͖��G��[�ad�{�)QJ���I ��d�V�]�!���n�2/ZV������K/�dvq��18��6�\� �3D�y��ﭒг@R�bz�;
����	a�92HTb,̶vJ��Qr󏐵��ǞY&W\|LP�쑝���k8���T�?�}�����'�EU{q`�6N>xs������q�!�8v�@e��Ab����:o�ߒ�䌨;�Y-�AGΔyy@ޝ�Q��rQ[�<Σ�q!�3���(�W-��!3���"Db�˗/7n�~���D���G��)SU��N���~�%2lH��x�H��X}i��F+���*O@�Ϳ{M���i��g�Dod�^ϼ�N�_y��K%;;U���V�-I�NB�x#7�r۽o��M�2튋̼�1��<4���W����z�����a����Ӣ��IP���R��$�3j�s�q�ع�M��(";��w�5���1��s&ʇ�+T�M�|�=�6�䆟ɏ��K.��x饚;���o�+�z|���6K&�^�lV�k�1o�ae�)�����1�R~z�q�B���ei��?�#/,�Ȥ���80ٹ� kښ�"9���W�LQ��@������a���r������t�/��q0�]��u�WO��ɓMX�
�j����c�k�-�!~��������-?��L84K�A��(��={kdgY�d�<U�~�ʪ҃H3<<�^�g��e�A�O7���]��'d☞2����k���5����5����Hbz�Qm-X~�
�_���~ ;�����O�}p�Y�#�z�� o�U�e���s��e��s���B��!����6�*�.���a y���c.�����TVmZ!�%�ū�+}�9jȑ���� ݽ��i$e����Kzn~б螷��{����-�d�ƥ�֢�FcJ�/��3ɸ��m��H� �9Vr��s6�K�C����Stޕ�p�j�_W">�aه��)�����&\p���I��w�.��]Ch���hH��5o��o��0ZZu�f��p�sN�d�%�.��1��*蝘�Gz���~BH�ə72rɽ�:QrG��6GecD<�1gވ��y�b�~��!8q���®`G����x���!?D�TĘת�!;"rq�o�і� �yc�3os(��ɶ�����,Q�z<z=o������jYhP�����/���Ӎ�E�	~~��a)R�v���E����(q���^��� �|w`�d6R'h�[�*B�6�9������!>���3���o���  y֬Y&I�"DCT_~?��3C��_~�e�k|q-��{���>������<���Ki�A�cSe���ciA�x�bg��xꩧ��N$�p�Q��裏9�q�Fy�wė é�hb��8
C��;��c���ůApjR���7K�����p��/�ɲ���D;�7E�Q����^��J|j�7�oSF��!}����/�-/�چ��d�z%��(M���)��֔G8;էc=��c�H}S�|��"b��_r��Y�I	q��Ty|~��'5(�N>"KR������A���2���*�|��s{��Kf�7��U�9���	y\����Izr�؊Z���b|��+���D<u|�Y��,,1�fGI���N��u;k�9A�"�oR|����OvD�����+.�
�A���� ���Y�Z!ߜ��hۊ��Uef�����Se���^�j`�D�')�����^6�3��=vH�D��mv��\T/[����2@L�Щ���;����ʥN�N��}�y�N��t���Qį�V#��$^��6��������17��=L���k+�̱p��),k�:�����|y��r���ʱ�3ewY�4�[��D�����d����g�HB��7.5|�-Z-�,t2�T-���|;fJ��i�qf�r:�Z�1��}�RX��K@liu���b䎹%R]��w�V P ���c!pM��KG�׉���qeO�yڮ7d��-�+�T:�_���JaSd��dx^�<��^5�[�`��v��� �����)HX��u;k���c9A��� ����<�v,�\e��x���;K䝏ˍV��/'�9�^�Wf�a[EM�k_���%�D�n�wV���"�Kuek�(c�`��݂��sXЁ���,�3�$O�VR٨�ϰ"V��χ�~����nWM�N��0&S��y�҈�rK���ݶeo��M���f�F�o�,��Ň���O4i�6ށ7��؃0�X �6,-
�@�HeQ�Zv�a"��.�!�Peez$H�Z�ŕM��R)�j�0 ;��:/,n��}q�>٧c㾌;_u��=�g0ySii2x�`ٽk�,��m�)�ѠN5��gL�8o�*�^_Q�\H��=��A��פ��}a�HGE.���ms��	b�ymy�!x[c�X춋��Dbˬ}�D�����t��ҩ ??_vn�&K� �A�u��1��'�Hz�7��dm�]'��WF�q���c᰽c�
 E�,t�
b�]�z�!�������-Y�dI����s�1��t<QE���铝 /-��� PO�'G������w�����~wbY�<�B��p��4�����	��������5t�Eň#�����)�h4��?hA��x���Z�I���Q���F�N����ފ�#GP�H��[��t��T*�\x�&�Ǉ�E���_��C�Ô��q��E���)=Ϳ�T~���)Ƶ�9 �;i��4)S�m�����~���:*C��
� ���Ͱ+`Q�k�_z�%�e!�����,N��ɥ�^z�����T?��F����k+Je�jZ�(˸ٱ�Z� ���6��țE�dD�d�^�a,��D˲�������׾&�<�1;(4� �Un �$\�_ a�wךh��w�E슺�f��o6!QU��d�aCᮓ�6W��?�Q#���F�ފƮ���$�m�ԩ&Q���g�}V^{�5C�0�C�������8bH�	}���Mmz����V�I��ũI>��iʆ>X[a��l6Ao5 14�-J/��U[��;�m��� �J�޽{��ˍ>����4�>EV{�]���o\'9i�&"�Ya����A�a��_W;y��FTq°tc��7u���� {�Du����!�	'�`�`v�]�$p�� <���{�VY�&h�oeC�BeƤ�Fi@y���ii�.��B Mz �%�<�Z�*�P_A��A�����e��bΕ�P���������p0Z/o�ʛ[��<��kd���6Y9�,�E� w��/� 6 ��&���o��8Ot�kdA�,�Tm*sd��4)��aCh^�J5�c;'�Xe�ʭ5]j��b$U�Р��H
.{�A�zx��ϝ �bx^rH�Y�\�E��l��=tGʝ�4�U6D���I_௯,�)�g��66ICWʐ@�������3�qKM��?�|���,+V�~G�xx�	D��xB��q�/�P)o�Ժ�]��į�@Ö�u2�"��+��x;�z�+wrb�a���W\a�	���'��~��"�����J ka�s�8n���W��eJ�W��H�����yb?V�w��&��������#yJ�:��r�9Bl�8�!h�C�&|�nۮ��pH��SO=%4�a�!*A@.>({�UWy\�=�9�m1(��x+�A-�uҨ���+6ε�a/GI3�E8��8ix��O6A�-E��dO�!R4�C�����VXTѵZ��#���$^d	�N�������V�ߜ�D3f�0:5�0J�8�7��_C$W>/����T�;4Sm�����Ę�qy��p�z�if�%H�� d�'7���:�Ⱦ�f��ۘ�߻:/�P]�~�_�n|Ʊ.�&x��G���r�6Y`�jS����G�L�/5����$&����� KA��1z�"-Z�
G��;��T%J/բrt�3_a�"sW����~9�2�_����u4v����+��X�:;�o߾f�����i��v�te��5��v��`V�*\�XIZ�Wv�8�`&K��Dg<�jXRhB?4U�	�l��7���j��
l/i0�t蛪��jv��Bm���׿6��/���}�٦0�̰�o��4}��H9bB]���#z��o��b�X�P� b[F���S�e��Ϫ�C)D�<�'K�&��OV{�n�z��ޙ	����bR�
.uv��nM��I�g��|C��j�W���Թج���׿�e���v�i��B���QG%O?�t�	`���`U�$�b4͇��Ak�l��3X��d��&_������l�ߐr��#6E�Ly�G6=�N���~]�]�Kl�&�Yw��	P��!�C5��&b2ā�ݸ���y.���Ξ���,Аȟ��C,��!ҕ�Z�Y��C|n�CM��RGf��6� 	v�8���Ů�,rT[3Z���O����t�R�ԅ%�ǧB�v�DC 8qb����:a��r���,-�=�fţ1���0��`m�0��cL��d��GC(�� ��"�q���թ@�8G�?���r�uי������T/êº:�C��
���O7�%���af{���`2d @T�'�1dՃ�}��mU����O�el7ۢ�g��tY��p[���SM���|`ކ�]bm�zWc��b��`:��7�鮩�
���������m>.+�,D��hP�T��)kPA�J��v���#�EL�ú�dk�ݠ���[���v�,��+�m�(+((0JS�XY��ّ������{g���a'~Za�%���U[�=���j#kI�ț��V�1��p�WWB�l�r�{�����$�6�j����Im�u�=XS��E�z�hCMK�aSM��C��@�	lu׉���k��ӛ����x=��=jQ7 ��x:�[w�6_yp(Z1��	p4v�mj6�W�.��'O7V�b�I|q_"�'�����&>`,�i�B���iӦ���~!KȘ�-f����9�,�]���h���� ���y�xĿE˒�������w<넁8��w		t��w6��-�Ƹl�m-+���&����T�v,��]��] -�^cx��e����i4�g�ظ0��}&?����,�lMp�E�����F�W>�L�vZ��΅��.M�ˌ�n�y���Hqe��+�ND��c�>����}Yx<��ᮤP�`����m�56BC�dkjM]`�4L���� ;X�''���J\�<�JEVzs��ek�]���B���D7�K!$���3�L�O"�c��H�ƽ�lm'#q��d�*��,ͱ�!�7,����	�9pRw�pX<oر�.�}�!dH@&�w���z<�|�ȅwה�5Y�!������RS��a���\��0�.�<ei����.�/9o��K�/�$�{�P���4&x�ǂV:�!G�H{Ƣq��.!��{m�_�I!� i�x{�����n��p��`�I�t������ԟ�����$�ט�	�o��¿��`ߤ�m�����E�Ŝn$�PI�h�Ð���%)�qR�
PA(\�+�և8'�H0;���$�C�~xW!���2d.B��¶b�V !|�&E��>�������� ��XI�����C�����o����>:S�\P,q.����lA�Ӄ7��X�ZSx,�R�w�{�9I��V�Ww�#�����BXԨ�,z
v�$��w�$������]l�F1l��-D��LS�X�Dd�2'V���Ǫ�k��;k����'c��I<c�;������~�9D���5�6w��Pv &y衇̿�Xz4���<�yYT6��Wl�1�8�:t�|[92� C�ߴ�0v��Ϧ�'Ȋ���M.�g���Tn:�B��?&~ī��P/��îx����N�,`[!�݀��7��w)E����1�4P�+?2E`{q��V�k:9d�U�_[Q�dǻ�b��|-�f$�� �S�F>�Ġ����f��զdAc�˟e�� mX^��d�����.&��O����|o�Q�ρƌ-S���QwESk��n�#C'���Z2≭�0B�o� �$����k�4��x��w�I�c�G��`�;���R��-m��Ml�D��_�u���pv��:+�DY��
���"���h��:��v����������� ��u[�P��@nG�u%X�XW;�ŉ��x��fnl=_[t�=�6���l�. ��8a���Z�C�䴁g<�wSM���l#zsP΋��`�0L@*�M"�z��
2
Wms�O|����A�;���
r�P� �]���%���	V;�(^V�0L[�X���ɟ��'�$G˾�
����o6�YQ���j]�:����,蟓h�������^|e�-�}g��dD_��Ѝ�������JJ�z�}YV��\d�8��sx.��7��Ұ����~����\�gN�a�uV�W�\]n¸Ѻ_��N�|����f{M���;&��,V?�E����vc!���j7Q�=�����o�&y�^(AL��D�)�yn��R�~��=eцJY��ڴw�uB�W��Ū�� �WB㯊�%`��*~9���i��<�m�s��`S�_~�! �qd,��?��pm)V8ķ�e�9O����������:"K�_W�+��$���J0)A�+�X	QB�`�B�:*9���f�,��)��b�R����#�Mׇ�n�[��|�?��O�;��E(�`q������t�����R��g���cOd�����،Z���C6�ݽ��=TV-W[�*��}��D6;��d/Z-�*?�<0<� ����;T~yzaI���_Hn�(�nvRLA6V=����-���AHV<,���u��֭w5X_�o� ��c�1,ş��e�������'�:�EJY�J:��^��Vk�(M6�G��B�2��S"���� �2L���r8lZ~�.���~� �����w�qH>/� Ų6��|��̙3M�
q���7&?�	7�tSTyb�NrA/,�ՂgFXP�s��qJ����%��#�#�ߑT�����Gf�U�+�7Jr�	(I��%��v���!;�`�P�ЮP����?���L�ܝJ�*Lw���p iu�4bqr�DZ�-`y�[�a�õO8,���+��-��>IF��;�p'Ũ;hXoji0���x��z������`Kz����TиPy	\a�>�q(�/�����ch�A	 ��Z�D;��aD.q�ʭ����h0�!ׅ��?���^{�r���{┅�G40�l#�V�uCa����E@��� ��|�»#E4����
{��z�3�zDT�L���J2(�z���`;`��4�[*r��⻂�c���M��n��CU���8�Bk$����b^��:���z�T��[a� ��L�	�/:Б�� ��K%p��!+��HU�_��2 ��!q�����u�����!��C���i)��w�)�AI��\�3I�q�v���I�&9��h2W
�;݃�CwH�dAr=2��*$X��U`;ʡY��G�>��!������ �d~����"��[Kq���x:�Vo4)�MF�#�Q�I���=g��4+�a\���z
�J��(�tw�sw����fL�PB��G�駟JqQ���^'�a�+�Z��m����~6!��+`��+���o;;�]A(�gzp)���np�Y�29܆; �0)u#���P��kdO�Y��Y��*�b��7A��7�4�����r2����<]3cL���-�����o�����M2�n(sx�����3UgD�#A��X�$~�Z��H�:ݼ�1�0�L���	�$����.uH�)vH��5F���D9�= ٰ)� ���ļ�n1l� ��d3����߲i���47��Vt��c���pD҈�ҍU!Z�7Д̨�^'N�)*k0��`��w֔��v��N���v�!m�	�����闕�0Dj[��rt���;�=���pʑٲdcU�1\ t����-��&Y�&�3_W�+ٚ�E�(ma��6iҤ��B��
� =)@ H�0����n4��`Y�nք���&;�E�����O���Nt�O�"�.�	fB��K�`��IT2���w^0Sc���t��t��-�u��K�J�k�"�	E�g�u�>$<��Nkw֚RU��!Ć@Se�T ��^�:�N���;��|�ȁ4l�R����f�qh�x�E���1/z�V����ɼ4� �V���0�9�͜��e1���6x�(c75���cu��7E��B��9�F�H�!�$<P�jGյ��!���n���������=���Bڏ�3�˻���\[~C�u�RW�}Rp�p0;{�ؘ���i�iJ��h�!��.`�3�kk	��t������ç����������?Op�G�6�ڲ�X8�E;��S�ۉy��sQB;�� ��[�����ilj}��RR�Ȥy�����벮d����Om�\[��VbFgǒ�F��X��JQ��,"�L|�qm!x5�$�KCRRR�^�DO�T����'��r0��Ma���w�3�y��k�KQѮ�;����l3v��n�3����W_-Y�Y��ܹQ�Hj=�~�"��?�P��|�56+;K.��"s?�T�_�|��m������7�a�<l��n��D���Jq�[O����9��2���*[\ �b�)E�DxVO*ՁiJ�F�y[NN�T��Ew&�JZZ�uw-�7��ǻ�yw�;��n������ӷ��y�Y&��M����7jēE2$?_�y�9���/͑x �X[�y�̙m�Yބ��hԿoU�?���[%*�&8����Y`�w�!+����(׭7K,vɐz=�Dmm�|ec�&L��OG��A$�G�p��	�| cC�h�� ����x�� I��v|B|̱�L<)QbE��=

Z����>�r�s����}uʔ)�_}�U�k���)���AN�Ȉ�
�ڮ\�T}� ���Z�J<F�]x���|9!�r@q�/E~�4ü뮻�:]W�lYү_�Dr|6�DiP�<r��1 ��C�@S��J�B�)}��:P��ލ��ڇI7��~o��������L|^c�������<�a��(Q�Z�飼����u>��]��������q���j%H���>��?m�,��񇑛d���J�A,��:.-���uXEQm�@�䣧���i~Z����t��ȓ�L��4�o���L6M4��L=�p
�yْ%R��H��k(!�B zø���j��`���^�'e��z�=d-���%�j9<i.] �c��c��l��p��ז:p�v�9�����c��Y�<(7��"[�6\z��6oR�۲cG�Z�>b����a��ٺO��k
��L"GF�3��5k�.��8����}�ň7|���6x����{�rsH �M��U��'�b �?$d��(��\��O"{���N��'�"��߼�̂bAd�� D��o�86(�����bR�k3H���hK<0	h������f{�M����L����?_����h�����s衇>AT�7I�<�0D��曏�gK�(Rv��:CU����SSS_��� ��I�2o#��DA4��JҘ��~���7�
�A@������a�}�"�.�}B���� =B�O���l�~b�7�t��7��A�%��6���x.�3�-[��3f܊������.**���c��`^;��IЭ��^��:�c�٣ǲ�s����۷oϡg ڃ�E &q1�R�~�l��ްo�D�Õ�g�,�Y�f�����E�O�0��)�'�	�#��Bj/���XA^��:���[шY�j] ��g�x�\�E�\嘚�(q�����ڍ��T�w�����>~�a�����n�՝oP��	�:0U���"���^��ICYE��lKX�;c�>����<^[ K�=���3�!|�q���ܰ.x0Z	�x�qӥo�L�x�֭�`ڥ߻\�u~��{�9�d5����e�`��W]e
1�O�S2��P&M�l�s����:|�OԶI�{O5����ȸ�ɾ��ED���1c��{�>37����S����N,Q�fԇ��6���@�=	�S��֣U,l��`_��
?묳̃�7�Y՚�.�f��#��;��ew.fơM��Z4��-��m�b�y�7�P&Ƽ mlm��a_[�w��X����^����� G��>3�S�e=��S�>m!Da�^�ν�xFp�BR�'!�8»U��X�p�Lȃ�'uoyV%+���ʰ�`�Æh�ikYm�$n��p  �@2Id��؍n���Jq$���������ޛe��ܯ
�q����]�=Hp�柬~[�a�"c1��n$�k�FN� A6���^�wV��31��@�� '�m��9��]�| ��j��f���ժ�zN���w7����hv�U�16>p�B��&��}^o`�/0v�~�u���h8툽��� �u�嚶ȳoR�����[�B�t�uy�1ʧ����Tu��3Ϥ�؏^|�ŧ��8�t�6�f���c���o��\��+���cC
�u���=��L��e:�P�|��7����M��`��f$�8�U��� ���3�x���u�H��={v��D!�x��Ǔ ���ĩ����(!c�{T=�V��y%z���_�W�}г�}W�ࢋ.�")Ĺ�+ڃ&���UbD�E0G���� �`�灻/��_A��A�|E�n_���W�f�A�|E�n_����[�V�Ax    IEND�B`�PK   ���XG�~��  � /   images/0739a1b1-a163-452a-a325-ab452d55b136.png�y8�m?�r�J�M!*IY��Ie�^Y&������[�d�cb�0��d�1̒,�ٲ�L������������|�|�4}��>�r}��|��mn$�_l��mۄ�o^�ܶM�i۶]&{w-�����A���{����� ��n�m�&�I����em4�6�l����
�*y�����x(����WŶm;����5��9t4Gb&��Ȳѹ�}��OܜΉSٱ������b��MT�}�L�1HƸD���?j��i͘�ǰf�	�A��{�ξ�[_����J�z���r���٢w��/5a��t�I��ե�EnhǶ-?����'m�ں-��Ǔ[�n�-��v<����xN��J�h���e3��2������7��=V��)u!";G?�� ��<�|K0�yY���I2,���^)�Ϭ���Ev�p�����������d���4���dK;!-�L�^�$Cx�䐦W��k��E���9謗	* P��ϕ�����S�����0C���~�?��$Ǖ���φ%mXJ����{���w/�y|
�T!��;��G����쳄�[�����⩧�U�6}3���6��{�[$��ab1�P��~z�3������Y�q(�V�f��¦�&	�� ��l.Z��s9�2SH�W�ơP6�[��SnT�QokF!s�Ǔ`��� 6rl�������fI�:�v�K�|l��%����)�m����}gw0�6=y�dk��?�/������<�w�}l��جJ���s�+����������6����Í�͍{3�����"R-33�	a\yoU+����̡-�߶~�S���v�ѯ�f��nY7�߼�K�pE߬�����f�J�\t���+"D�,�����AGf�H��X��i���&���oց���A{10�^���l����UL&0���ٵ?���E�)�Q�5��s�=[�,�8�v�Y����>\��>\+sS�N��88y��</�!-Ot�HS�/'9��q�ZwuR��
���ӝ�v�����xS>edf5�Ի`��Z��/�j�3�QM�/
�1Q �wH����G�h�p���"[�|���fi�h.��-
��f�:�[<?>gh8)�2d����q���j�GZl��Ϩ�4.{��F���Hq���5�1͸�m2�2~�l����]I���J�&k�-�x�T�/�O�z�5�k����8��JdX��a9�<��V��\�����R��9�����0�TƦ%r�hm�[o���b�Pԓ��YپQ5Y�� �>[Զ�f�UG~����bhA�A	���6��,-��:[��Y����p���m���k���A��p�ʂ�K��&�{sdJ;?=3�O�	}�Ij�>>wE�Ws20NJ]=X�uq�g�j����bN���|�G����Q�s˪�r���W��ӕ������7�[����v�ЂF�K^��FY�{��s��ʻ��R�:i��D{��x�����T�Dr��j�M�s3�����:u˙��[�.�[Im}�v8��0��d�Y�S�ܷ�BW�V�F��V�E��V�
���355;����҈�RW&/�+�'��]W�e����v�@$�Y��=�Vܲܽ��ٳ�6�tinb��[s!ޞ�C����<_��iG�Gn���_a+*�� ]>��-u��{\lrǹ��x�|�b�ߕ��?e��@�㕸�����[�`J�p-��i��m�'���n��:l�xm�pd�l�em,W0Q�:��"�A�fXDyP��pOTG^uPiN��c��+l����~ŭdyώ�ȂrZ�����?���A�Xc|O���/�Pc���>���tx/��g�N8^xai=���
\�ΟNXi��@�l��]Q�0��!a�+ץ���q�����`Vq,�o"�B8a�i���Itq�����1C�06�J��J���
�<-VTy�����kQ
�ɍ������p�F����Ϝ����r�}��O��u�~�Ar�u�����Wc~2�ƪ����@�m�����
&�H�;7��.2g�>)l!�(�|�v�z��[�TJ�й��#�J�:F���R���:oȼ�>33�w��vå"����P|�?{�&��#�H��+���#��<o��Jڐ(-�������&�Mt^��R��|٢����q`�g��c��j��02���)����F�;W������+�xR��:P��/�ސc�H���\k�Ý�/���d�����^� u �Ƚ���c��������-6yK�.�d�j��܉�x�������7�.{��"�'�>����K�۰o�g����m%���UY�> �/��
zo��X{_�v��Kû��q��Ŧ�ү2#G�_Z&�k3��x��r��2#zל���@�[��װ��^_�L�#/=lql�X4Xm������nq�p�7ME]�A��J60��e��ogU.Ė�FՄ�W_Ћ�[cT���l�hze< &��x����/{�"�Lv��
��= з$:��Ln�_�|_�!��ɬK{U���G��Jak�6����������R3Ć��S�ۿE$��|��ӝ1��E}��q[s<w�R��.�$����V�P���Lկ�0e�YK�9��qO_L���p��Tu��/8�ˊ��Z��]��A�@(�^�1���s�z��'�l��x�}u��A���<�� m������j��1õ��B��iB��	�A&q��6�t���+�cQ"M	��յN�I/&�'9�˹��Vv�t�R��FAD�/��"������N��+�',��Z.����xT�;(a��C��?����Drɴ��J@a��m�e��h?-����b	���M8=�^����=�ӽ�b/��Y:#�3���rp`��$G7��0_��s�N���vo���B��
]\�R�	�e�1cٝ)z)A���۹����E;DO�V$���t+˾C��@;�sA����.���8yQ\��Gwz�O/9s>u��ř����e�5o��e=���qפkx�t������]�o�O��V��f(�\z/�x�@P�p8��R��fU�j�nL�`v\�\fM����qY�cGr�?�������@�W����:��7[�zȏ����{�N�ND�v�bKT�
{���=��s,�{B-#+�Vx�Z�%��/�(?��9&s4]���5���3\>�P(y
�6*���+����&�sN}wT�$�8���/Aa�ԥ5i[����x@�� �`��������4�nc��,��R���1��q��a��­��[C���	�~n���7a�F��G�S̻1[�#ݹ rŀ�}�uNʂj*�6I�VU˕��UP�����h�1G�2�Rs���Ծ�y[�J�梵3d������A���i(Β�����~\@?�,�8�(ݙ"�i��ݤ�܇^��g�ms*$��ESפ�#-
!���U	�����lQ�̵��K�1u)�ױ~Q ���16������	���8@qY�&C��.:!�6��;c0߷s� ��g��"HSK�P
��10ڂ�|���}��([��`�d>�*��I6�c)<���H[Y�ғ���,~ �lvЧ%	Y�m�[��>+�8U�t�@�e@��v�AB�a������m����p��_ \�**�>j۪��q�E'|���s��}��)��Һ���w,���n�b*� M���1?VPg�>V{���M�|j�:`�@�������x��Ox6���Q���s5��I�a��P��'��C��ݽ��(��/(���Y�<x�̶H|�d��kѺ>�Y�G`���*"�r��l��$-.���A@<��E��u�#�n�����,�=�bB�B��^ͧځ[�<C��^� ��|�C$S+��G���.Ԟ�*��� AP�	�oe���W�\t ��i����� �D=CZ7��<���?��1����m!�����;ZЮ��|�-����;����ٱ��rO"���_�yF�
�`��!�;��U��X���t��(�JW9�~�#&�M���j�n �I=�x)��s�Y��rvHYF|>zBf�؉P�":�m��'(����n�?0 �捻Dr��Ox@{٭�Qh�BU��_FQ��(p��
�zk6=U�E��+��2p����v�)��Y��4`�n}��Ƕ��.E�Tes��q�e� p3I�k	Y�պ��ľ̫�}�Q�@�i���u��<��mЭ�6�e@x~_�"^X��$Ԥ����txY��&��_�/薳�q�1:z�3#9�Sd��V������#�����m8./����V+}����� ��jm�*~Ԉ`*P�,��\aK ������=}�������1�c,��s��E��J��3�2doR0�e��&��}
�)@h��}�G,;�`�͉BJ�Q��ib�]M%�%ᖝ�$�3���0f����9��.����l�O�u+6��,w\μ���� j";+k�Q@��7�HDi;w��d�N�Ž�͊�BX���+z���I��Ӎ�R��2��q�:�r��Ť ꛕ�4�J�\Dt��>w&�����Q�)�,m�k�b��	�KM�PA9A����C�T}�v�٥M���dҊ-"�Ҧ�^���o"�.��Jf���Q�^#��B6��&���(t�f�4��g~yŪ�Y5����A�Epq�3���Ĕ'�Д��*�AT:Vb��|���-%�uw�e�I��UU<��2Pl�SF�׋���t���ޝCɶ]+�7���Ld=>e�_�T{�+�F^Tx'M����DE�o�-l���P�G>���Ѐ]
�?�8a\I��$��B�Aِ�"�n��P�j�����Oy��eDH��t�k#�AX_�&��O�-���T`g��JK�7J��"�Ÿ�(64U��]'�YP��D���я���rZ~�xy���uu$|�2���d~���a�sa�w/���������&���5#k��'+��}PkH,h�d��v���Tϴz��Z��G�_ZN�ad$	c���Tx�4�nʤ��6�P�����ʞ���|�uxP�[�+l��VF�߃)��k�~1s��Q��"���c&�,�Ƶ�ͦ�X���ϠoC��l�I�v�$Fc�I��2!cY����RI����-䋴X�Za+K�k��Z��\�=�Y����n4a��gT���SQM����܁G�"�]������ ��wl�q-��/\y�u��f�ň7'�
�l6:�9��#�!X�Ě��b�����F����w�:N[h�[�n���=��C1;����M9"〧����;/Quu������� ��N�ۖ^$b����|7���V�Â��a��s�.X[�H��M�K/�evTv>�U۟��gSǄ�E�|���Hr2���}U{9��y,{�hh����y� h9��&5�Pg��X�s2� �b��ͼ�tzer��;�4O�+NfpE/�ݔ��(BW��r���9����(�oB6������픴Lq�K���xRtJ�?K((2�~^>��npM��Y��#�)a��ݡ"�#�|�a�*�*�j���[e�G(>�D/��(�|y�W^ x�m#�]���h��0T[fLL�j�~Ԅ�jo�u��9���p���r~��So��}�'�ť5^LP�1��
IJ�p�C2�����IJWC&� ���/��\���=%ݰ�){�����{8�ގIR�v
�Hp*Mi֪�X;����SAe���x$��V+<�$���s��\~�z�}x_a{�x{���#2'ͳRl"�/=?�z`��V��s����8�>�ȷ��k��*98��е��zy�i��S�h�4�?_�\;���Yմ%�V%��b?�����ܕɪq�ꑝLO�t���RT�^d.��p�*�> '����'b�CU/$mް�Q�ql�[�3@��pu��ToV�@���Wz$�jIgg.��]bT��$%
�?�H��4(eh��Խd�,�m��cn��B��
�b�9�uLT3��	yX��a�*O��;۬&����Ⱥ�6Kо�S��`�\�˙o�
��Z�d���%�����隲��/�@,���z��҈��I��cW��f�HЈc���h�|���Z#��Rt�Kj��N�\%�����n{(�ډ<��3�r��AI��֞��C����Gz�.Zm���J\i/��I��)�k|�c����l3	]݄K����'�q#��+��?_v}c�1N(��ߡ��~5�(5�T�Ӥ�O�!��n���0{HMWǥ<�����e��ؘ298���i���|IT�VDb�*y�>w����$�Om�~W�z�n�W(���r�
�z��Kȯ���'�q?Z�X���U/7���3c�n���e�����հ���e��Ym����� DQ� &5��}z)t�ȩԻK����k<�q<�2�1���<79��������8��в��u�F�'Z{r��(ഏ�,5O�o�ܙ�v�ʨ���Sn)ړ	h:ͽRj����D��j<s���Y�H�5R��z=�B���㼌��a�}���UZ�6�@d5�b��	��sV��5�n��7n�:�m��!�'u�	l��1*�Pte�
(���l��U��<$u�{�<l��F@�O���Wyl�@�+,�)����a�
e��k���O�X3��J{n6�Z���G�6o\�]ʚ>��R�,�g.����{Y��ma
/0���U�υWcnI�*%\��W�+�V�`õ�x�����b"�r�=�\����Kmk�)3��g3���	Y{�D�}<�76+7Ŭ柕� o�|feQFW�C�:?��\lS������[7tُ`@?����چ���� }zY��E=	)?YQQ��-ח�q��syBk�S�3Q�0�w����`�ӷ��FI�e�c�B�g�Y���_���x��l� ������l�MҦd� v��q�P�>@_�����^ZiE>�)>���K=��*�ڍI�t/��.%S�B@�����T ��/��GJ�{�fm^ͥy8��ro�Vö�ϿNo����i���ѓ׹F4�6�>jY�::�zֈ�K8�Ϩ]U5�SX��k�<����)�Q_���ߙ�%���sY���}�Q��*��4f�d�Q��*VE�z�5�
xI##:@�t�}��+�{�;��$Mr�J�������/�\��1x��U1y(¦}]ĤwD~���C���ڣ�1��H{�g�d��4=�Qa���M��QZ���ը��fGR�}�\��8Ғ�q��}�4;l��/LoF#�T��7����֍1�ޣ���'-�xT�C��h*��-'�I��M�ڈ�s��/�_�{�����G��L��z�����,�+����F*�޳V�����>S���D�Rg����;�m�.V<�����3�t�`#����N������M1��nܩ�7��u&�]�{جʦXO�k�௛:Rg�L2�4�Z��O�TS���q֟[� ���]�h���uj����X|��Vmwa�O��D�����K6}���n�Z��Oe��b�u��2��A�:vq��L�J�� C"<��Z��������������;��X���H���[���jB?�ݧ�#��Lr
���-T:�+�D֗��@�E�ѣģ�|Qgp=��F�uK�ܫN���Q��� B���Ƽe{\[7ҵ��H���n5֎6�~�b�.bצ�!�P�	�	G���k�눸������J�|������^B�^�Y�n����5��f]$g�(M,���D�h�t`&ȍ�f�j�7���xYg]�22X_7�����=��f��7*qKn�ֱhUr�Y�}$U��G�e��_~�T�1�;��j&�>��!��I�.�*۬�=��(��0T�	�GU�Weh�7bTQ=5�8�n��މh�\�_����+D��YZ�wr��V1Mw^im�G��@S�ɚ��� �w\E���Y�wStH���n�
H����v�.�ѥ�n�]Ux��D^����ї��ox�%��!�����NKx�#��:LۧYf<�0�W�z�4	ռ\agM�*�L��2�^caJˊ�:������Z�&���DS�zu`;%4��P���f�e�`�c�wH}�*6@v;���9_�ġ%�]���gƷF���S�T��0��o����� =^=�
���"�����P8� �ױ+^���#�3*d��T`� A���F�>�o�{�҅W=���ʾ�3�yq�z\�S�Ѩt����):/���G�*����fZ�5q^�3���XRg��X?��p�O����7p*�̄\���-��d[�P	M(�vQ���nS8�Z���j� 4!�f���&N!���[>��^������c���
��Er����ֻ����۠����q�c�]G�1}WUv仓!TE��d�*u��㴧����ag�1�Qz���,���R��yI�u�(֫�^�6_kk���	h<�"��Dk�y���'�ߋ�n�)�k�K�ngX,�h�{�]5Q{�q%��:�Dв��^ndH�P�m�R��
�>lB�D"�tf�����^O3�e�z�stX�g%����u�	��<�W<��m�Y� CDhkX�� ���fß�| An�G
�H��`�h"���L,���;/sC����HL��/�2mnM�� ��G2y�d�of��;���>$�����m=SfM;��&��n;	�,ů�)�Nl�]��3잡�.[;;˦��Ť��Φ=w�^��i^���`�#I������X$���}���L���l��4
��~Ti0�l8 z�Qٚ�(�~�y��H�`i2�>a�S��U.+׸��L��TO��<��u�@����#	�m�s��ӆ�u��*���~��fj�6���>�H+��m�8�B�������l==F���t��'Y����eo���|��$��tT
n���W�k#e��ND�\nB��.�l�,���=K?����p�|[��5��O �x5�L��z�L��Z˹H������ׁ�3�F�Q�Mr���4�4���2k���m)��4e0�$KufN���'W������L��3��̡���i��t��nQ�eJ-�X*\p.22�	`^c�9ν�z,p���ş Ɉn�}# 9|z!D�!J��W+�g(̏���\w��>�����	�O1���.��p���׹��\�h�(6�3��d'�jMk�XC�ݺKc�E���$K8s�1����m0�# �
�Cln�#z��gI@�gAЅ�t���:�g0��Z�2���	�1�6/L��%���I�(.-�}�g�
�)ޔ��}��_���OrV�^���xK(��Fe���^��"6�w9=��1�k�k/s�bQ�1L1ԃ<�)�N������uac?�{kQ���>��
@������R��m+q��j0ߕԓ���	&�Л�軣����b[`�����\�:��s	��G
�� q��H����r4K�;@��]	�D�Ӹ��$�����?�	W.@���)������%Eg��G&�Z�ɫv!%�h~�=p���~xjX��(�߲^0k����W��/	��kмj��P�
ʑ��Sv	�E��1~��R�)+L�
Y�� �P��E������=���WH�zq��{�3:k#� 
<.���?O��H�v���܍�M"r�I�c(��A�5�Ŕ����،�z٣�B5��~��tI��t��X�}�|N7pf���M�ڷ<fțP^�̙\}&�"׏L�p5
x�R�1yQBxV���v�T�%+�������j�n�	��E����#�}�z�-��S��G�=qN���P��76��2y�ɚ�����pQ�XW���4 ȤhS2P��+ZK��s؝ڛ��o�'���g����l~�`�f8)���>��z�����V��������?O��4��o��A�ΐ��&�d������^$�0��ٍ�47.V����9��B��OKH��<*S�����Gy�VJ��Eu8������\����)���kYp�<�l������'��|ݻ�NA~�ֿidC�量s�Tiy�E��r��x�?>W�F����N6a^����}̶Kn��
��-�����>��ݑ�O���ܡ~��3� �(��p85C���pR�n�{D*�Y�`e���zb�1�L���a�Z&�AE|�/Q�%н��]�d'�� �Vx���X����9ݵ/��t���n}"���%c�^�����u#}tD����@OK�IT���͛S�&��#7E�bή��>����գ�$?�o.��Y����DYP1Ёt��#��d �	�F�7�o�vؙ�s�5DZ��[ �w/�E�j�A�y����xR˚���cGe�����rO�I��d���r`�#��7�<Ʀ*Rv-:vE�ُ���?[��N�l�`0��_�����/�����4`0�Rp��3T�z*[�'�L�:��{e�]���z�	��*���I����ފ�j7b��~�_	���8�)��PV�z����D��8����Wdg1|�z� �(�߂]uB�p�:�%��dS8���Q�B?WE9Tt��̀	�ǋ�v��7��,Ö���ip@���ڷ��U�s�}sk���c���;���r�>l ʾ�����K2����"\ف�{>�!3 E���o�.����7��D��vv;��Zu�b�&(��_��eD�>2�H�TA�E#��s�"FhAb@j��%Bm�@�Yz��X��'hN2>��������M]����>�T����.��ʂ�`���<!`B�ju��`5r���`"��$	˔����T�F@�m�\�(k|����;c�XS�D*�}{�!ODC!�x1W`G����a�DG�z��B0�;�]�!� �q�F����?�8K�I��0͠����0�C�0\{�>�'@\�Cȕ��P?z]�*�1���e��C>@2e_���(U$���#S<0N,�t��i�;������'z��'�]�cDm
D��#+R���_Պ�����a^�����J9�
S��%t�p�������9�{�F�N�ǂ��;=�?����_E����g�Z=��;��4�2 ��)��\~����"36�(��C� G�)��T�pN�s��*?O�͂�rd�Л�_&Ϣ�{���vX�v@�;Iϻ�^��tP�����p�?�CG������+�D���o�s~����~ߩ�Y0�4��  Kn	�T ~} T��a��u��J��}Wn���NRVՓ�v��#]��9ʂd]�,Z���̭L Ț ������E��,�/�DM�/}j��HI�O1��س��m����N+?v˶	o�LQ��6�W��@\e�p��uZ2+7�&�����~!OV3�\�Q�c�0۴9����wN]C=��%2�N�b�|��ׂx;����t�E��4L�+��j�d6�YO+n�YUMP���ɜdD�=`` TΙ$(I D�5��^8њR���d�e�ɰ�}v߸п`Q��?��{t�LF�/��k5�Y�#b������&� �iw
:S���\�Q�vQ�a�(��Ͻ.�%�X�z\]��J�K4��}��<�ư*9��isx����?{�㕙* �(��z�׸��Us��:^��]V3�M�߼?�g�皖���rS���jjS�s�g$�e_2'o�G$�����I�w^��'Ӻoh�"��^��W0��rK##��9;y����܅,I� E�ӴMa�sv�!��?�t��� jG�7ښvD��΅�����t����s¼�0�������f�t�7��(}8�"�>�����7��fTP�Y���ٲ����A�T�t�]۪�pq�఑$JF@�@m�M����]��P�7��}���˽S��@O�!�ҵ��n�׹̈́K��X&)G�m?a�S�U#ah%��	��(��+������Gyw4�L7�E�;�r�\1W�}������Rԉ؋����R͚C}Ύ<���:<�����q�\����	�d
+I�~y�<xxQc�F�&	1j�6J¾�8���,r�z�]�U\Уv��.<�M�]���6�����I��B0�a,�[-�����C�o�0�qcè�����t���m��y��`r����l;[��j�7����_�:�����°ԝh��l�k�^;�� c�eIv��9�~}x=a�{R!w&��ݒ��b��v��gO�����\��:ټ�?�[Zڱ�i�	$H����;�\3G�s�k��"h��]3�oz�&@�NV�	B(����s8�WuM���؀zw��(eJ?����,͎ø�o�����1/�ʙNك���A�]>?��bby�H�������OYjŝ�.~M($k*���AD����9.Mn�w��sۭ;��WJ�u3�j�o���� �8]�Z��Ͳ�`�:��� �1H~kȃ���h�g~ã �m{�xJ�}���f�;_^ܽ��<k��>m�&p�h�������1SEi.Jƚ� |N��0� �#�i���_e����{+/"4jS��O;>��g����rAlP������/>àÛ�Rʓ�`��r=����*�U���G4��_fx�"�Ǳ\�X�A�9۱n�5���1��kЎ��y�-��9�1t��&�=�����hN;�}�.~7o�qU�+��照E&�V8W;Ͻ>{PB��ދ�z&'�������	���t���LgO
�,�9?{����@��`�7��������!���[�ʔ��H-20f#!)�99R�4]���IQ�T��f?� �o�3��>�%X0{�}�R�2�GK�W�5�l`o�AK�4H/����dwh�>-�)��o�C��.�r�C�f�����^�b��,9Gc{,^�9���9�u3����o���&�����j������-�T����،�=���t��������`�T����=q�����bff^���@�ԧ�m������_�ܱĂ���H���vr������=�q	7�Rg����_I�/-����|؛�>uɯ��BQ�o����Eþ�e�����A�!�;<�uz*}�wa�N�����&wr��?ȟи^�v��`��ԺP��͂�OB.�,r���	�߲���q��9�?;�Hs1��s��#�U�Ӌ��*��2�o
�n綱� �7g��J�-��u@M�q����"��ׄ�v����Ղ���vW�T�$������S���N�:~k�m��Tr��X?M��nU����a(��̅��o��i@��[����pj�rNpX��W��?�h�2�2-���`�W��/��*����؜Ps
�8 �� @��ݙ_�c���5�FL����;qA>� �k<~�Y屼�G���ōv�Y�7\/䃧�F�J�8O��.�Ҭ�w�;^���ӥ���64_�����
�Ƨ�g�l�N�]9�z�N$Pn�v6 ��ƤK�@���PZ�N����fM�*!��}]��`v����

 �)!���2CJ�����L���Ӭ�>��뭠7���;����@��egXa�3��ay4�w��)��/|)u�4��3��]`c4��<Iٰ|ԩ��T��Z�#�l���q���^�������<r�3{���;"��
Mw�����k���L�j{���i1ڕC�ch�3J6[�#Y�
�o�i�f�u�Z-�@���|�.�g2��L>�	����ʰX������HreA_�pw��[&�����_�{�Wq��pL{��U�w"��RMk����2�zœN<��>�4,M�z�B���~"�_�z|
j�l�T��Q����?{4�����~N�_�ƢE�v��H���ϩ�#��GO��M�/�֑�k�.H�s�>\s5��I�&ڇX�̒��g�0���u]^;��d:�����S�K@�#L�{�od�F�,H���c�\1sZ)5���u}�{B����L�5�?�T#^�:G�-z�u=�ь�FG�C����s�u��j샱�'��|��{���C���|���<$11��];����#Ъ��]4;�V}s|�f#���|НS��� ��m�J(���t55��E��8���K�=�)N&�}���U(�ׯ���w��(����;�%�RWu��J�Ś�I��~��KA��;OV�@�~>���TI9�cz ��*@���򈌴(��	������{��Ps%�n�E��轶g�;*$P��U9��5���_����wU������޲��*�w߬�P�D"��f��"��\v���i��T�ſ�D����'л�?�?�c����������!��*�r��Z۶�+����8�W��N4K����0��P�=A�Id$u�ߪ�-�S�y���m[�aT�����Kw��x_�ȷ��j�������hg����=���������7�0�4�1����@48�Iix��<$���1I��gb`/�V��R�l%��'�H%F���m��=����[��=N�\|��(��	/K���J��γkpۆ��ew���&��r�1�Z2���@`������lbj��/v>��y\m�@�J�0�,!�r*o��)<���QqaaÝ@	r_˦K�d���$�����k��m�=7�8�a��.ľ��S/�F+d�d��]���_���9K�9�ڼ�KO��D��sh�����=}|e[�K9{U��햲>���v���8�O�ʥl�U[�Hx���$��Y�/\��Y�$N����F�	}}P�!���==2�:h~]����y��cQU�ք+�5����LE礮ŭ���
�&3���O�R��u���`HUE����;��:(2S0���1�|�Z�RTW�[8{0M*���+Aj?���!nm�4��&��9���CO�ZF�v���|��.�^�kz=����V�ϰi��=�։R7�|�!hR�� �Ra,�7��&՞Q˺��.��#�vg}����2��B"4C��/�̵4�}�QֻXل��%oj�@�������h'$ЪX:p�¸�wh��	���t�'/e.83}���<.�;���8�U�z�������"���==���ӳ�?Β�:+���=u���oS/������U-���?ǳ{�)9����:}VL5�)���^��.��Y2ri�g1~��em/�{�ȅ }ȉ\�����ޤ����� ]g[�M��޹ժ��q��$�)]����(������)���0��j֧�Q~֟Y����A�yוGEwThe1/�67z�ظ�H�J(�''H��t~Ş*���Ҹ�ϰL�̐���!U��"�Y��f���g -����2���j̞�(�p��0��]���v�z؏X\���̫�=.�jk?��[W�V��o��C})M2_x٘��-����|1�<��JU��''�y����h�P�W�#��������bvM��e�����ְ��2~��N� ��M��F��ͩt����ʼ���F���U��y�\Xp	�Q��uչ�0Z�*�nԔ��;�!�k_��CN��x�E����PM���<��i�AՓ�"
����E����������^��7-�e��ƙd9ʇ*��x��JcJs�>�ԕ��M=�EC?x�#\I�g��3U�{7&��f=�Vwh� �l\l�h��t��+��
8��l�e��h&���7�<���)�'�Kf	����ːDz�r-m�C*d�dl�ou���"(�bV��_���d�#��a�4�`��O��%�lӑ�:
)����X�B*���������RN��
��sƁ��� x�)�+�����.G;�G���q�_����F�(���G�~��>�~_&�6��0`��(�[�\�N݂]\����t�?����s7^���//��s2�PK3��� ����C�FC���K+]�)��GCi�H��tG
���&O�ݕ�bֽ�:^��6�R����$�Ԇ�Ig�g���Q�ˣ�j�W�OX��W<�����DX|�����Uu���qu�	k�Je�Xpӕ9��)�d8
�Q�a�9"=g&���A4��wL�|���g!W�<�fJ����oh@|��|��N�`w�;{�>�r-W��nN�	�M"�}i67���#Uvß���+����eI�~�]�3}�eC �ؤ�qc5�
Z�:�z@��5(.�Ƥ}k�Zs����J�?1�7k����<�����xf�	����^���$U��.�Ս�7���7��q�gV�g����t��Mgߛz���j����Q�?:��������;l���0�l)�J@�@X��'��jwx��پ1`��p����~|�<�	>R-��鞬G�M$�_x�i휱g�i�
�7$ cE��ɸ~�O�T�L�I���o_����´�nI�y�/$J�L��ȆA����2�׿�F�GF�=�I	��a�_r˟ ��P��j��3��q�iL�N�����$��/r�J�o|���~��bMuuC��E���%�[�*R�{�����ĭ����c���όI����K ����u:�45��i㫴x���CM����8V/�,1 F(sa����j}W�I�{ZH@ڃ�NL��zxA'9��p���PJ���`|ĩ�֒�h���CO����t
ujL��Y�7�a����6�����w�o�x�3R��J;���t��h E׸���z���7�KX'�x��ڢ�ULW������ipw���x�M����^]��;:E1�b3�6��t�'�OB[�0B_�i�6���,���Y.L��y�ܙ�F�ouZw��O,3$m�r�}��6�>Cx#��t��8�����QM/_ߨ�c��X�
�DzWi
�;��^#��HWz�{�� ��.%AZ(!�����9�G|����u׻�k=�יٳg�ޟ�e&|gB�/�!�>��	[�^l�I��۔��<$� ��rŒǅx
-V�-��T����T��h9�	��oXi�&��I"���yEH�;~�.k��b��MԊ.l��d���u]���m
��3�����8'	�Z�s^eh�����<9�hW�!j�S�w+GǪm����o���%��#*��x�������i�]Sr�ytfh<Y]�4��i?O�R�/h�7�$]��ث�f��\W�=?.-3Z�X��e�.5���'��8�o���7�zj�3_��g�E-S�a:k;�o�3]�Q�j�����������&�y�b�kJ�:%�h�R>��9�!j�+���� r�)��(�8}�S�۸np	�}-�hI� RT�L� ���<���fH��n����``դ�+�r��E1l<��
B���LrB����G��X�c�[Hd��<6�� �/o�M�R7.u�����qt�i��ǰs�3��\��h�#��ʇ�]�k��|~;�L��y`�0'�D#�L��J�""*��#r��6)�^!k
�����`O�Y�0�m�[����Z	>'�g���])7)I��\��6��*��8jO�SjB�6�ȨUW�m���Z�=��6-g��X4OK��K!i��@mx��=��:@����"r��CE��"��i23n��FƬH�S�U�Ca���m���Nc9R�i��,2�Rk�4>�y&���H��^�OR��cl;���*Z
��Y���\��&7�X�s�@��w���Yw�~ W�Wǵ:���E�B2�s������m��#��jz�}���rV)�|+I�յ�y� ���7&06�5}O�U��/�a�+�~�b�m_ �f'(��޵_i�OR\n�@`K��p����>�ACf�d�<�j�wgC�_���B�)��6�ͯ�ne N��_�FA�sRG�{ô��� >Qį����U��:s�zOp����551y����8́�����G�������.�k�5o&���(�Ɖ&dd���F+�q�=�Y�"L_�G"2,�T�嚡�'��ܵ���)p�`��p*o�C�EB|s>>���!}t�挿����qZ �\���mK�W�G)��|s�Ɨ����s��k��s_���d��#�B7�1�
lBR�EH�u
�|���ǝ�Qe���%�Ñ�u���J��%͸�4��O������~�"�͢����#0�OHK�ǃā�8�ǀ^�B!}S��F����Ȭ݈��j�ykG{�A�P㞣x
�o�USu�Q�[��ټ��!�
e�T7f�<bM�īvk��ZȦ׀�Ɇ�j�$2��N��&��ϛTCۻ��o�&�k/���u6���[,���6!�2BjK���x@�轅+�,;�2ʻ�n���úL��ب���:O�Yq���5��+]}�0�b>M�[��V5*VRɄ/���ARՈ��o	��<�v:|���`ϰ^Z�ƹ�I�C���ܝ�:�TY�$t�Qr)��}�jM��CTS�k���v�1�諸�[�b��nv�;VQ�resK]�\n�dG����'p�b�V�L����k��m��_���[n]4Wh�gGi8�"RW�h�n�ʷ�!���Ş�$�3�n�w�-��"'��4��o�	�YWB�H��#�3h�D��_�mA.���9̳%��q�Cb���{����Xrz<B��f!��E��[+tX�z�(P�rZ�`��z��*68���E�m�NY&����n��<a}�(�j��Od]KA�vN�>�e���+]�
s���'*vP+�>	�-�6
�[d[��Yj��oh�*�кT�:z;�38߲� ���ƒ�8k�vW�7g��[�7B%�c-���M�M,�*�q�L��.$��$�w�?���=a�Q���5)�$�
ۋҰڞ�}��s���lU���^Dg)Ќt�q���[��������)�&�>��K���6��FrY�`{|QU����=�20
 �*6>��$�O0=�U�Mbّ��L1%ios�<p��l���ot6�m���oI��V3b�xҠ���W��Ob����A未c�[��zq��8$�����:Ӭ��\�o��Bܠ�z'|���I��zẶ��[��5D�k��+��
�J�'W4�����yߚjYE�l�%6΂��{#��+�_#�{�?�9���X ��}�U���n>g��͕�x��C���Z�~�9��ۮ������DX;h7��wH���~�@@��d:t���@��%�P���i�Z�HLLY<su����u	�⮦1���}qa<o�x�9�e�?n_�|�RQ�
�gT�>�g9z����j)@m�T�V�]�l/&�~�r.�*�A�{#w�dլ|�:D��+��T\}!��³���#j��� `��:�$k�ڎ��>0$�<@s�[�9}q
�K5M��$�y���"�'�k�Z���E��M��|c��:��+w�e�@�a|�;l���V擖�:]X�b>TVw/�2{��)��5ta��U����.�k�3��w<���ٓ�ҜD�1$��σVk���k����-�{������#h��6�ŝ��LqVuSU�`kN{�嚰_�M�.��}�@}��ul���Li�S��g���5]�+�-��`YTu��x2.��e�̐hY2�~�=�j(���UU-�7�&|����Z�"[�%���dt��W%Me$��ɒg>|��U}Q���h��{�=�4G_��x%�1�w�^��R�Wy�[�̩h�h��B�[�B�U�r���Dҝ͞��V��-0"(vߍ��X|�����*���*�l�DS���d��Ed�L�[�~G;�f�Z-�ж�%�Ȁ�|�>�~�@��Lh彈��6z��Ͻ&	e��J� LOot�:x��Zg�Ϟ#��(#���.�Y�L[� kC�ի�.������|�륟���a5m^�:V��Q�T�c. ���X�	�BϹȂ�fe����99
/���YZ�h�c���Щ��A�ac�fӢ���ojA�_�b͏��������ߞ_ ��z��I���:/ r}�,��C "l!w,d�{q|��Ǟ�������sVα�m>�Z�D[�N�85�
�m<Q����)w�������C^EnQ�S�w2��X�D+��J��0�Ub� ���Ė�S��r!-f�X:m|×/��R9���7ƽ�4u���]�&�/i���Ѵ�>�`�rX��,�,����q�ߏ�����jk�4�������$S�t�Œ�����o@$�q-��L�`6�L��Aig���gc�ᶂ��p9f���:�����F�i��}|�.��E��+�ɴ��[}�!�377!V�W��v� ����(���fūj1��i!S��w�x�=x<)���!5����~U���)Db�[f�:S�i�4�+Ͱep[5MS-[f;�/-�4�S�mX�g���e�8��E�nIV�߶��<�IR�D�+��s�
H��ZU0���Q�㙹��%*�D�r����-���G���w�����׊h����a��-R�U ^z/�_-�]y�e�8;�M���+_S7B�4�
���Ro�y�m�+?	����\�ݫD*�_��&���NI)�;t��&yñ][+�"թ�!y��˙�z�Ֆ$YC���0�e��[|ح1ʽ�y��OM�zܭ��|q����VΦ{U�Ѻ�z��֘��XS��y�"|��;�i�x c&3�ڷ��k �Oi��[ׯ�6�m3=?�U4�ݴu��x��#1�x()=ׅ7��'��B� ���Y��idr`�X�oH����5�2��=K�hla�h�l��MY�^��$�N������Y����*�� �R+����-;��ؕ����kƱ��[9���{o�XV(����P0O~����NV c����r��S�E��"�6���@����w��Z݁�#"]�b���)�(RazG-�UC��gp]�9%�dw�r^)6tt��pҷ� �7��uX��g)k�5��q�x��G�
���6����^K���x��0�c�sQ�&�H����a'�7{R;���l?��X/����
Q�^*ik�����8a^s<e�" ��N��-�9�t��u��!P-�����'�CAէ�W&�r�+��f��]�߇%&a�k>���>֯�����JW���U��Io�� ��^�������޺�ni�o��t�_T�u7-����C�$�H�l�7w`�k����Q0 S�[�f��~��I�\��Q��'�6���L[͕6eE���*�#��	Q���3�R?ې�Q��"4[�3����ʘ�Z���eM"��\����.�4�\E��s;Q�i~�%X��X��@�G��?�9e#�~ �N�DV����X��&;a���L�)��6� b���w�9�����:��>z��w��7���C�5�&_@�	iI۪�|���F=��lG�2R޾�wyJˑ�{{�̱O�_U�S$z�3�O�qЫ���{���E*#1�x���P$G����GƄ� 5�M�'�<��|����9�SLf)�Dn.@K�׬�D7o�Љ_��6`6�^w Չ�� �2�+� �D4��(�^�m������@�᯼E�'��C�șq��d�Ze����D��]�.�+����:�t��ʐ�5�>�M�w;+'v�pX�<9O�������r-nst�o�Ho�P�����ֿ�<�H�LW��Z�eN2��4���O����ؕ?�{?�id���;�9t5|�0��M����'!�O~���ᰣ�	����E�>����)c
KV�z=��v�cv4Qm�]�%l{_�/���J�z�DԲ%�������T:�G�� ǂ��-�k�=p
�h*_.cr)���b���n��B�����M����ŝ�@7wT�
�*�u}��ļ�>�Hnd�m-��t�S˔`��mX���?'[ǭA�64�3Q�E��u8Έ~t5xխk-h�3��	���f>�9�r��i���t�m�W��x(��;N��&���C�ig�L�K�yeMHJ�7+<��T�I�������U���o�,���[U���@l{�zh_+��~��y\T{�Z|
AA��S$:w��	!�YUa�|�u��C�^U�Ms�����Z�Pqc9c��V�/�a)�
�~�F<|'�6%�jk�)��@��v��x����6�E��EK��+�rx��u|PH�	Qq򉶵�{�T����O�ԽOڵ\pL�Ś�%��S}��pKqE����'	U��8VP�s0��\:�T��5�(<��'�K�Ι���5.�������"��U\��H��"N>X2��f�p
[�e9� OF��4�(ܴ��ͼ���)��t2a���(��R]��*�
�2y B�0�,�
�I/�{_/��bsw�y���??~�U[a%�3`+��կ�DU��ǧ����>��1Q\��
�l�����<#u桅'�G��3�������@��:�[��Q���a��N��м}�Ĺ�*���&W,���.�8Җ|�t����%U�Bk;ij��gpM�̅�v!)�\o�g*���bm#I����a������P�!;�X��Qvn3OU�L<;���tENe�[�@fv�p �%��s=yd��ѥ�~��]�]ҹ��N��k<YZ��Tl��c1���1e���\@YL�Pop�R �[� *�솆C�XS"��R�O'� +?/��$���U����N�z詡����-�Ƀ�-������y�z ��`o w�ne����~s�>���2��Д����R��+K�M��]��tų�Ӽ�%(ķ,a���5)n>5ޣˡM���	>��4���;��N���R���2��R��&�b`�\� r,s�����e�$��D2�ɑ���jUG���{i���XOmu��[���T܋�3V��%_ҝJ^�:K�2�����ƻٳ�P;\�~ϔG�)�Н �|���R�����m��r��[W꼟�Fi���ɯ�6�|�^�^ee�Ʈ�trL~'�݀���ee؉)e%�X�����u{}N��:�!��l�4��n�c���b�܉m�?��CN֖̂Qq�?��@�^>�f�&�ȃ�[o��M�B��M�"xj�O���l�=�������ǣո��x
�iǩ8��|��s���׶8iw��L|_u\�����c�"��il�1�>?�*5O6O�@�����H%r��M|P�6n;o���-8�BK%_	I=~܋�ۂ@HSVAeU�LV�򛊷�y��t���=ҫ� ;_p^y�T)|Y-ϻ����\4!>��z�B.�|��҅�<3{z��Psv��Y[�Ϗ� �L�6b'b��:ې�싮�,����=���7�$��,'�1w$ׅ����C��6
@�9�J���F%Bt]u�*�+���4�#@��߿t��*0�iZ��!a��I�VjOc�т�qq�K|9��'�Q.4Wڐp�~���D��9�I�)�y��N�
Iic��  �A!��n I�p�`�p��[q��9���6�HV��`�WF|	AVMw��/��H� �QTJ@�˶+�Zt��5�f׾�y����8	;`��H|���a�zk����'ʧ처�S�v �Z?fIﭠ�1��k� �X!��e����^c(D����ߊ�y�E�A������F���)%*J�H~DR����K�I�,ѢU��A��;a���j�]��-� �0��6�%���YEb=xk��5�Bt�h�$��R C9���N�����ҧ���&Egc�)��7�:�(uaU/(=�H)<�ꂊl�\^����L�D��JS�G*!��Թ����6�U��O63T�����R�W��NIt�z�sڱk�`0�-3	 N�1y�S����3�"�꽡Bg�B><4�d{�$	+b�Xez���zԞ$@�	K��2���9�:\d^_�݃"�u,Օ��n�UV��Rd9��s`6w9[�� g�?l���R��c� �h���cB�b�������^��*�q��9N���*vLZ�������e"	�أ��Kޱ��$Ia*g%��.��9���mXj���/�1�j��@p��d�f񑈂�dʗ�X�S:�l�.f�w�e�u2�߾�dr�}�<(��1���k�}��sJ�Xm�̩J�.��`�GGr�ԉ��@����]3��������^LG�e��O�2G�n�"�� �7��aʬ�ry��7�ۼ��}b!�����Ĕ��e7�WW�Uq{�H9)�ޤ����O�b�G�x�T-�gK�'Bh%j�2��>i�����ȴ�cJ�/De0[3���c���p��'����ȳ�N��&���%H�o���3s�u4)9}|�=�*�,qV����߲{�+�[���_�L��XGY����d�m�nz�ƽ��%U��2�Yʹ���c%$��Y"������C�=�`���Hy��*�C���@���s*R��CDÉ���Д4��� ��9|�)��׿'I�.���/�g�}1���������,����j������ ������~������I����w^b�����^����?#���S�Bw`�������86�L�C���0����^���%���|q���9=d�4�+�ލ�l��!��]�dϮ�Y��5�:���-����%@@f[�J��'����@`�Z4o�k8gԋO��>�F��$_Uy��D����L���o�soߤ)Qˍ�1k�T*���Qd~����'��<����c&%>�:�=*�k�-�2[V�z�>�f^���4}'Xh%�3���Ĺg�X��~�~0J��d���po޶�ŉF&)�CZ�&�'H��JP}�<��f�*'ihV�����w���D�2����}����C�AA���Z��U���{�3��߭2f_�N����7P#:\�`�[�Z�ïa�8�}�+� ڟ�*��Y?���pMv_)��2�Gz5Ri6��t���:v1^�^D��lk��Z��$Iվ�WJ�܌�v^K��%li����~\�x㓈�v���(�!�8���w;�E�&�T�������
����Z�+���^��s�c�z�A�Zk���[UM{�����{�a~U}	�g�0|���RH��^��� A�|$�x�*�Aά�����"vW�n}#��r$Q����@v�&�4�[{���Y�غL����M`���Q$�|xq�xR���#l��#J6nf���̪�J����7�V��g{"���@��}�-|*�&	��|�y��
8����s6�����e2%��
����X��C��}�U{�T��
khO��
1���C����9�p��
^����:ع4O(�mJ�A��g���!���{���+�M3��fP�w�&�OG?�|E{Y(B5\m�l[��'��l����Zo�ը��
�����aJâ��K�M&5�-,��H���md���<�j||>"�>_�T�r����~Iq����[�}��Hy�(TM&�`��i��rGn�t����,/2R��!c�V���{��{��۲N�ǈ�@6p��&���z�F߷ �=���!i������S�c�2!��C�%Ȃ��;z�b��c@6X�=�j�ve8����4i�2sF�೩����(��"C�À����a���`�����pn�NV�H�p��C�FDD�33Ծ���h��AO��+��e�&���ѓ�)��|ȉ�B�rOxC?��D�����9@��햎ײ6��c'��y(9�a�v�hV�黎�X4d�j�;�����+�v�T�����8�#Q��d<���õ���-��C��&���cD\D��O2�����+�`��J�VP@�́��Z��!��6�juu���>-GkX.&ᙑ��0�hw�¼TRp��W �W���u{
,>MaB$i�R;2rr�Za岦HUϖ� 6r���-Y�tH�;+�e!�������wH�@��P��|V#kV�ݬrO&1���8�ٺ�Iص��$���?���o�lg�I��D>d"���L����hM�b�(˚{
���ha�\Z4\{�*4�@n����k��i�o.���8	[�t<��q�(C�6"��T[$��$�d�~6<��RL�(��Ob��)��\ �J�]CB9��e���n��,��4Rqp�b����gٿ���T�=C���i��{�l	�Qv?��Ņ�W��r_�C5��;�K��V4���0�ј�[�﷏�=�[�٪�����ǻ�Ʋ�~=y�]�9-]ћ��f��f�i�̺!�	�b�E�����(w햾�w�Oy�_iٵjﾹ;)���}|��8jt�Qvɦ-� �����OD�����gt�m���'�䞻����!'ݭ��ok���W��Z�N��}k�L|k6' ϻ��~�����銿P?v<j�J����?k��vtH���J��x��*D���E��.r_+^�����D���+���$��[f�;SvW����J����t���5�����U.j�	' �nw"6�@�����0�W���,�+>
2��씎E������	���QI���0��>�ik�N,��U#���p��r�p�ũ�V�}����o�������� 'q����,����6�kLW'rx��e�>'Q�u��j�����S֛��������a �7��
�t�Y#>��#�5}Oj!غ����ݨ*�*%8�U@Yp�έ�njg�ԝW���a�q1QG{/�-0'D��������/�������L�/�V7=^�{:��R����v�cJ�h|���\G�,���SSo��*��Y���d}���iX����wT��&�0��M����� ��U���jq�6eA�����|�H���B����� ������!<.���@\�j-$��%�^�9�M᫴/T ���ơ��;�}Z�Eҋ�V�9Mm��և��ߤ������TdDT����i�0��9�(�U���YH\p�f�ïL�<��,�����NU�1�bg�>�!�7�W��8~[��!҅���<o����}O��А�]�������i'����:=2��m�^�=�E���4;��z=W����t}���B��#��%Mb+��k|ޡ���	��@�PuZ�l�ע+Wv�y\�eWf0���:u�i��b*p�}={|2$ry�2_�ʊ��7���5��1��&�ۯ�����uK;���|5�=y��4�5x�B��]T��y�(B~TOA8��6���$N�p�ˬj@ZyvHh��jrM(b���i�>����(���-kr�TŖ�����u��Ğ��*��z}��k�6� ]	K�~Ř��p������=�.O(��~�[��Z�����\Ӣ/́��/�ii��yը����O��%�[A?�H�>��䞿N�%�8&�IW��ү~m�Sǁ/���ܤz��qG�Y�,Y�n��ք�zD�!�����e>+P��vʫ�~�=������T_�e�>��|�wJ�"��z`�T�+�;Ojգk<ޱ&�]o�Ђ싮&Z�2Y����D���)j6��p,*��֏�|(�@���E�?��M_�[ �*\����缋��zE
N6���s)1��6J�6�������rDG,���x��Y�Jջ��iЂ��B�|n�E����2��4,�iN�Ep�݌ii���T1҅T`���]���W *����oUS����ʆ`��<X����3 Xx�b�@�!�7�\����!�!�4��3T��hF�Չ�bx��M�}���i�K��+��
���<i⦛I6NCwz��m�v�F#�R�r��5����y}ҥ���7��N`�*��½���s�O���3Z{7+-��8��ֆ�V��Y��7<�i^��;�4eP�a�hi2�2���ᕧ���~J���<O��%�Q����%M`�ƣ'��9c��)�.Þ��Z�*NÞӒ���g�6D��z殍�:;b3�ӊ������n�e�秫����\N�`�9��������<v7���Ƈ�$~o�y���ޢ�:�0g�y�%0�w�Ea��9�^伛��a,�M���;���P�T�)�3l�%���q�>�S�߽ݱ�������]��'�?�)�g26�7���`���D<+.��ۏ�?��L����)���DN3�����79��<�ʜ��%�pjʤuֵ����	=�n}����M�S>�O5'���k�1v�[Ke�vkS�.�����ݺ�)(,l�1�����h�5',q\�MgX!U@�Ĭ���5(��{m���W����9uSS�A��������k�r	X���A>�<+�U@��tБ��=���̵Y�WB[͛�$<K����EL?ui]̺Ӝr-f����w|��*��>W'V5?>%��c�F����LR�u��4ۍTa;Af���G���*��n:�R¹/�|���8������[`u��$�-���,�������ӞZ�0_���� �RH����sԲ<�<���GaR@��y��+	�Wn�?�ʜ����%h�!��(�l.O~��Z��=�*�DI�]:�S�G�`���Nd��������kVb�&gm� ����'Y=�hO{Ƽ��}���N�X���
�����[�\�����?t}�V�M�0C���o�\'�>�P�?��d�Qʨ����1�y�[�)G���j�n��8jf���z&�Q�ityr#�Ϯ;@��IׇV���\�|ˉ
�|!�$"BWɱ.׆(Y�Y;+/�x������^���z2�U9�V;��m͸ں���Z��+�Y��8��>��-T\^��T��Џ�䝒cq��R��m�\�/�5a[]��m,lEJ��Y�Э�4�9�ǲ���c(����_Y��[�d����B�}v{�x�f��?���Q�������r��FW����䙩��r��`8�礭��kK
=��t'x���-�p���Q'</�+))Io��N���O�b��A/]����j'l>�^s����Jٔ�hy�ONӽ�g����ya�f��A�C����'<�.�� �Eq茈���O�/ӎ���%i���63�����e�c�~}o�>ͩ__���i&F<���W��i�;��ӽ��J�u}�6��Ox�衉L�n}���>Gu��(g�ޝ��[�O�D73�jڇ�����?��L9l`N�~���@�J���Ldtt�#�^)��� ���`ϵ��G����՘A�{~�]i����z{��3ix�U<1ES#{Ү��Օz�E�i$G�׉j��5��ΏlG��� ���QZ���B�]�Q}�~��Դ]4bc��X�s�����JK)X�y�ݑ4ϬfEۈh���Z� k�iJ0��6+J�~��I9�3�1����)������E��(�ds!F���pv�쌘5���^���y˹��4V@��f�b��#\�~mmm�di.��$E��/��;i~dH�'���kЍ�&��K`0��Ȅ��$v`T9������iJ�w���]nz��?�9�iv}�c_D#�#��� �:�����N�>���L��c8���Xdd�ܑe>�<k���MrV������P�;�݇�9z��`�Vs�P*�ƳcQ��=;;޾�5�y�.�;9bؔs�ڵkĦ)^>>#E£iJ���-����BQ)�T��Shcy����]�X�&L8��M����P�@�k�#��������QUMmֳ�d컿�q�<1������5S_jSߍ�_���@��5���1��!�6+�MS^�!�V����f�L$f�/uf��)�n�a��]�_`5ݹ��3�4P���:&s��۞$�#�7;e��t�5��\���gmy5�5k��$Tf"�C�'ݺ/�w�^\�|j����K��5-�*R�@�7ä#n,J�����p�NJ��� (l �!�TU	w�^7�t�KH`��l�%9��_?;#�+ ?6��N��g�Nv����u4����e�d ����uj#t�jCG�l
]hQ�A��陘�\io>0�244�Ƹ�O����t��ׇ�\�Ħ53X���1���dB��8c�O3��,�ç M���K�����0B@�!��R�GA��۪|Ǧ�� ��T��$�۲�w�G&� @Q�m�!D��N�.�y�Λv:���`0M۵��ݑ������@+��6�e�7f�SRRz�R�(�Gp���L䔖���!��e���?��F������FH<�i�|�y��n�%�,/�.�y��1C�-kdj�/x�HR�ABH+q2�;��}]A�f��<�:_���jW�/s 	hӯ�B߾���<ӛ,�ׇ?و>�ݞ@�_E�n���^�1����E4탊t
�O9�`�m�h4xm0n��]q�{�`聑��z穆`��mf8X��w����!t�;ݦk�w5�1?7�K��������"�[�SJuL���#�c4f��C���0W@� u��y�ޞ��Q~%�X9�!�~��+°�gv�k8T��y��<�"�i��xe��z����i~��>)""bfq�������ג$���`������?��������Z�ciP�a�-jj��s����Hg�b�e�8��4�d�FW��ו��Wk
��.N֗���</�{7���B��<�#[��wt���r�4�Hp�~oy��Yb��)\s Ja����a�!��K'�!�F!��ԿkN5��5��f9�~���fW�A�B����;�q��4��#���5�%��y�ɺ���ݼۍ������,.l��m����Gwc.ǜ�>J|� ����̧O�0U=����NN �0ź��Ͱ�wu��n��������i�����\j�+�9?���ܻ��.o�P�>|k��33\�~��S#kQ#���ܝ����@��XǫS��aL�!��g�ai��U4B�	��e�c>l�1|I�N�X����7�1}!�ߩ��s�{�������xえ��ʭ@w��&��-H�w����[I���΁?����.��~���j~9�k�_�\/�:�Fs Q�#{l���3���.����us��=dJ���J��á��GVN�WjD����"��O�?ן
=�ރ�0�a(P
Ŭ�f4�72u��F��4�,s6oJ�(�j�� G\�%աV$5�cI�'�;�� �#��A��i1�[_Hc��G�N�`6�N�W�68���!�� [�q[��Ą[� U0���s�Y﮻3��̑�3^ 7X8�:|bpp0P��� `�����fA̛f��/.��{_G�����:��*ۀRpv������	O/��A"1t�]��JO�ز]��׵�k#�#]�ă��*�@f��� �6�0��U�u�FĕK���~7����y��0`��r�գ�-��uu�&N���l�T���B����>bȄ;����*�s7���s�K-�#�K}H���V3E�B�w�q2�1��o�\��^�4:qFu�R�̐V��iAd2���%�.|p���S��[�}����AT��Lp�]�#!��5*��pM��Xp����#�rt�$���Z5~��>�	w�e���C�B>�(y�i���|�ږ�C��ߵ?y��[�D�`�(5�"��i;ފ��̯�@j6��i��V
��_鵌�Z�o�d�{W�<~���E�#h�l��$�\jTS�8ɥ���Lpв/����s�QGBنPQ�EA��7!�����k�ZD�+B-�f�c`޸��t�"o�T����'T#8>�F�
����W8S�����([U�F 8J������k<�o'�n`�����3��kߍV4B�Y鎬��ݻ�o��A��7��N�T-�F6���g��PB.;�*��J9�+r�/��yF����X��8���zn�T���G<�QA�a���ܩ�a��^��,��
v��/��sFiՇH���s��>�q�'+l�J|�1�d������B�xvv�DyVPa�R�e�0���6m���M]<uȱ4J�c���X���ɽ�eUs�dnGAv����p�� �R����9E��z����fEw�W�@��.�1� !6I��b!�HH�R����5.h��K�0;���1�wO�"À0����N�s&�1��5�F]�Y��Ai,�Xƨ���2�ʉZd�&F;{^���}iuv�{s�3Fri�?r0rf��$H[�0ȌX�D+O�;�B{��#�6[3�x����V:�@�Vz� ��:��X0�r��2��'��
˄*{Њf�x��	O�gb�N���O�t���7^~f��B�|���l��o����D�*�R����l��/�gEWk$��r� t�OL��˭�9����i�w\jN�\ҫPS�4�*��6y�`��CM?ɛi,B%$� ��j���oȥf�@���x3���#�;�Ԝ0�A-�.A'#f�VWW�b+���m& pU)�rt���f�I5�yp�<@r����� P�O[m�un�D��v����$�Ù����v�����*�I���f- H��v�Gieq�(�xfZ�8��ˠE��w?�a��0�������/�������C������xV���X���R)oeH�D���>�7�D�ĿI �f�������B�P�_��kte����
(��M ˰���#<ѵO���Ȉ)
~ix��7�]�]��a=�p��������ֶ8�wx��r���QGy���/S��	eh���TR�_���,��@��@�u��31a��~Y}���'p�w�^�����`C3ޕ�~gL�swt�%5�H3gۦ"��2����܎G��.�|��?�.��`�/�A,I[�z�4��eʯ1�+�s����8WY�Ɵ���IE������	�i��+�R��p�6y���N�Ǌ97�Šo9����!<I4bsrA��+h]k:
��5K��J�L�S����:�y|�PF���O?�mɓ�X����_�'���yY�/�mG*� ���$�d�T�p��d4��?(�%�nx,��)�+)� �o�G��d�F�E����;��[�*#���s�L�~.�%���lu}eBr3�>�t�n�h�z�pt��Ȧb�vK8N�`�2<��F��3���eƺK�d�te����6?�س����{�G�7��e i��x�r��椄��Q��$(��P�}>IS���%�'����� 	A��Ί'R�q��3G�`϶5N�bHT"�	��PWJ��A�/�RM��G����EN������
ZX�X�^�i�_ڒ��`�s�\U� ��Dg����B���3�&��&�0�+c�v��\BQ�v�`|���Y3�_�4�ܴ:�s��]��/��iǀ���|^瀚���)p3�!����_�T����_��_2Pל��z�+��?A�_�����s���1j@��?~�e}!j�B�GG��$��?Ww�O���i����E:������6}�:�ԔRO�޺����ڰY$Q�8W͘)���J;s��٢��SCr��z�h*G��@��������V����{q�j�.,��ڤ��࠺G*�j���[�>��ͭ,�V��&#��C����)�;Cھ�OteJ[���D�C�#�#I�LD~����������w���Sh���ƛ���d]kh��
�׈���F�֫�5:?���&�4���&�E�ѕ���W�]1g�hҢ���}�-�(3�#�kلL��`H�U�ss$��yh6�j��[J�~ֵ	9V�[���f�O�'�O��K���eX��Z.��ҒJn�_ɤ��aF�8C��M��@��4� �n���7��}]�]����$4S;h����Eú��]�5��_JF+�90��r�:r�͚:���s�Ṕ�T���
�l�j��}v2�ݻK����\3 9"4�u�ɝ�\:E~s$Ƨ�}P�>��K]�������2�,�+̻�a�S�ow�rG$O[^q��_0�t�|��k��ނ���'1w�'�row��H:�f{M�U:W�ƅ�"'w�;H�֜���7vp�mR�S%bg�y���J�;�rJ�y�'��6&�]�:�{�ѧi��{D��azU�Z �yb�ۃ�:����'C�[�8~ћv�Unx�Nϣ۠c��_w��s�=/��r
7���gs.����PMfQ��#��)�FP�)�;
�(D��4�HE�A:""-(ꠔP(]�H'�z �$�������]�w_����Y�q��s�>���v���\lUu��n����p�e��^�i�kWJn�b��4-��/z:����{�y���hK���q&�j��|�{G����e@5���mR���ni�q"n?~pb+��cV
4��� ���58�w�����Tg�ON�-@nn�Ȕpt�hB2�>Ι��^�m�c:���f��n�x kr��6��M��{��n.���]��	�^��;����w4������(����?�D��O�?�D��O����Q,w�}��t��������G*�a�j��8��ess3������.S>�.�6��E �M5;ח�fw��<G}����
,�KD�r�䕏(V�M]wi:��Qz˽�w�ƈ[��N�}�<��HS��ȃ$�Ra����
@:e�I.����x���pj��E.����͔p�4(ES,w�5>5S���_��Q��թ.��:�q�d����*�]�O��_���(��.��k��B=�!���|U��5B(��t�X���n9,�U�P�0��f�O���Fn��g�WW%����{��}n����W¹��~��O�
K�����=>����V^<�${�n�۷o��~5�T�P��RI-��um���dP��k��9c�4qM�;y��^H�/^��@��gyp��2��Í�Ύ��ן����.���<��}a��dT�_�)/]�F�r��)D��oom�ඬBH��<QUES ��HҾ���k �=��q����;Z��j�[m�;F�����	e�=��%-�g��V@yG��*�_�П"���'��FH	���\�t�α�[�Ł�2���<K���w���~���'kO�	��Úl�p������Y{T��2tJ���H������\$!g�7v���1�����#�#45��^��@�!�j�5ߏ�Z��A��0z�֤�hȔ`��LW����`���!Ͽ�0O��No0�65���]L��X�ʽ�&?���ի��mi�j�,� ޣ���D�%ni�H�!��r�cD�`4)A�љ�<��n�����3�a7l��(pUY��u�8��"qi9��bBi;m���IF֖�J�?�)�:�G�G�r ��sjϏ.�˯΅���\��2A�i� �咱��&�=����DG���1��_�V�yɸh�;�<D�x��y����It�����0�#��xM,_D�*t)�f�K7op}�%�q���a����m:6|
��1
����
�?z��Z���!G��l�y��,��b+><q���@\}D /}��~4���1:\ӟ�}��h��?rZ)��u��4g�����u)Z_M�zN��; �E~>-qͪ0�>u^X�M�M���Z�l�%&�ż^[��lME�Ѫ��PNvRMJ#�F*[ :#'Kp�?��yq���l��g���$4�1�fu̪��*������N����T�ՠ�'�k���u2�د����[#����jl6��p��+���u�ܕ�A��Q��oȺ���E��L�����?o��JQ�BQ�ZG�
�[�UK�]S��#2���H�����x<�.�8�5d]��{���
�zN
�覻o�����\*0pjE�}�@v��}c R?W��w-�p��v��8pbǥ�};�����������_��y�����/�<k��!��`-���Y�l��dԗT�������{�\�דN׾���6Ɂ����YJ�vk?>HG��sg �0yQn��k�4F$�5Į�b�Gx��U u$H�>�]�k��`�<�c�b/o�D]�^�����7f���������1?(|�:�N2����1��wא��{'جn4��>R�:��#�<f���L*|ϒ5�x@V��Q�k/%4�
�
�uF���'�$��n��A缢zE$T���������f�\C|���P�Θ��#��RY��819���I�<���o��C�XǼAZh��+���Lq��M#,�X�8N� �4p&N}}������-�m��c��+X{A�������>�=�F-����kLh3��X!�����m{�p�{jf���c�����y�BE�f�#E\L�L����+K-Ǝ,< {n�0�Cz;��\y�L����M��2�����:����Ck��}N����������TmJ��h����u�W6���߻܈���1��E{qa��X�z�*35�	 � ��C���}��E�jʜ7�z�LhC"���kGN?�x�&'��+�C��ܷq�/`���
�������y�J�W�@��EB�_�#�&S�����?����
�1F����ӉK����"�&8�S�[uB�b
�T�2C]+�I��ty����,��@�x,@̺��7.5v�/��>* �/%.�>�V�^w�J�#�x)�����S%[|�/��;�o~� ?.�,��&>|�l3��t���Y��������w*�=E���� #��sI�ƽ��FD)9�k�B:���IS�ݻB�]C�W6��;�_����x��r��y+�I�0���ɩ���o���|Ȑ�F�]��
գp,��Yn�u2r�ע�à����K����z��R�,�tEҾ)����{��؍���6�X� �G�G1um%$L��I�j����e�0�X[Kv~�>��w:p�z���ar���p=�L2:��ݶ�풏X�d�q���]�#*\.�#�ݪ�+_+�2�30�r�j�������<G.�~���
oBյ�]+Ei�׶2:�z�!y�P�����k��]���t�A�TI�����\)o�{@\�F~����2��_�k�^%��(v�_�n|�-O���H�Mhs�z��Iv��}q�k ���mÞ�	�]���@�؛����,�w�Q�qKaa��X*�R��<:�J�S�`�W�iK���B	�C9�,��������D��'� h�o�TI!/X���M���5z�ڷ�/�Y�qĕ��\�C^�����������ג��$S�ʹ3ل#V��r�O�ؖ�p�w�f�t��}W��S�\�+�7\�N5���f�]�p�"[T�D��ۏ�_��uvv�f������_�.���{�a���W����>�5�"�KZ~���J��\S����^�zspГtGW�� 7;�#xq��7XM� �i��D�F��u+�{��|����[����{��Pp��J�����Z�?��=���4)���a�hz��GD	?ݺP��	-�VO/d*wM@M����
<fBU����eW�IYɺC�1u��S��������5���H�X2y�5V�@޾�+�. l�5�aeƄ[n5aM4�Ɠo���S�q����|�ˉ
�(Ș�����K�Ԉ��� ���/�	�v�+bkF�Q��#?*�Ԟ��vШ�~��|�����xA��R�~�T�^/oQ�0e�����Ƹ��������\�91��A�No��?�bR?]Į��)&&�%���e�U��ѽ��3�2���$�}1�DQ���[��6Å3!	9�o�6�?x�T��G��e`�Y�-+,999_�\G�͕"��.���܁\ȷ�X���\���Jy������Gp��L_;��y88�䎳 n�����*K[��+/S�_���3n�)�K��H�[���?r���u�#���<V�k��s���2�(����B�Vl4U��dqa�3�
f��ʄ�X�$;�',�����yxr�RdY�54�D�>����ׄ����O4ϑ�m�G��"��ɗ���P��}C�Q��sؔ¹
l����A��'ob�pw�>A�q�7��{�8
�hi���8A���=�d���~���$�Y6̄Y���e�^0g��}�-�˸R�ޑ��m	���8g�4�ח�ó�h�3������>7��>�o�9CS��5T�j繐G�B��\�3ԝ�����`�}M�e#�.�vK���*�]�������u8>F������e]ԿC��u�O�L4�.��H�*�nޠE{�F�uӏ�E2W�
/�+X�	R]��K�)�B���W����u�?����7�ӝqoI<��v{�e+�'�x�VU��{�h����=��:�eQWV��R�bg��vѾ�Uh'�n-\�Q�/m�
���&]f*P����8.(�����d��:3��	!��â�;����7X��>r�~Tu�=gb�Z-�>_�["H�n/�a���K�{<`��,:o�;��ci�V`�,�h*�i�XU�g���^�T�bsr(V�D�����U�_p���K��ÂABe����f�:���q�?�V@��RQ�L`na�ix@�Z��ܞ�����g���.Kp����Eb����]+kd�vz�����,�>�;�I����p,��Ç���]k%��$Q}}}���:�5��9�E�������r���Q�t-{䉵d��x0���>x�<K��3v�����0��m�� �����y��䃔��&뢗�'�����i~F9!�UH	4�Cu�1�� g�濖�L��؁��Xy�r�\a�V�Llnn���t��S�N�-l���'hӷ
�� �;���/����!����_�	N
F�zf�����dt�cFA5���^�UfA�Zu�9)i�lA�d���WTo�	z$ ��F��P���n��|�����B`�N����G�Xg�dLyy"�>�wB��߇��\PX�)z���2kH�E��Ӧ�;��#�:���t}�6����5��Kd�����}��X�L`��.��~��P��&=NPY�N�n�,��/�|���S/��g�/ʮ�vyX���]{b�滆��3T�d=<�$�Xr?��CF����gryX�ԙ��i�����*��0��e��\;"�ps;j�jr}Hr��%�6����x�P@����i��=�]��pK[��[J2�R> 0�7�BKl�/��/
�K_��	��t��C�LNNc�c���q��=Q�󆼞��^0��Oy��Vg������ e�^,N�����d����.+j/h�Nq�6�U�&���Z�fbr���`�>�&��lsFe9�X����[����5)����Q#�|h̢+� z=i���3.Z�<11QǔȨ?�4�� me�p�IS��
S���Y ��".`��ԙ��\��ҏv��_l\\���n<;P�Ԕ-�Mt٠S��(�������շ���`N͆�_������q#F%4?�:UFU������rz�]���~��\�[M�n�g���>`�S[[[��;�����Ph�67w��7�39�-���
���CX�3��yh�R��j��H�tvvf�'��X4�<`Jj����H�?�+F����^;pr�����e�I�+<]+ �	�zzzZh�t�B]���@�%SiQY`ٲN�\��R&'ݔ?h����:]�V� mu٢�f�&sh)�fK{�=<��P��-ҐM���N�@�~s�5����qxju�K��h��lv�2L�Y�ͨC���{�3��
9��S ��(�7���_�+oI%�b**-�X��(ⶵ٩I�#\e��d��u�(]PQQ���KNO�+@00�Ծd��|�UN��DGGG��V��.�����)���n�,Z��e�nL|�tG�e��fuH�����8���>`)\�کEq�F�E?�����Ō��f��i��"_���(5��׆<M�u��b�B3���<�C�j}�x���އM,��:r/YF�\"��"E���=�v����|b����R�=�W�ta�޶�璋7z[��~�y�Zٛ=H�^�C�o��)��s���=3]���_w$�;o2p�8������wށ8����GyR;@���v�ꏷ�99�������/�Uȳ��>������y222+3]=��'`���*�����CCC��&�}��:wy�?���9���������_h��K��P6��&ݴ��ٓ��̃��%c{�K"4�Z���4�~	B&���1rUN�h�td�#�GPs�MH�3�%�Lm�jӛcb ��q�t�����c��;��]�WٵJDPWV�+��.J=Ӆ?Z��N�3; �#��!��1N��iN+�TZ@����B�vu�-7������k����p�?�꯯�N��y���V���o�w����bS:7��Im�����M��D�����a�����_OA?*�<;��>�f�_��'?I�x;9�Ư��S�c�Ϝ�{7E����W\��h�	xv��ġ]��rq)Ĥ�9��t�`3G"E��$�����S�!�>�D	�%�B��|]sՇ�<����K���"���k���p1���� ��vK.v~�D���G�OS�ͪ��瑧��9�iԖ�Vw�,,縕Y���r������!o<_	õ<����+��������n�D��7�_#���NC��V��i��|�n�m��˜�6q�&����P���Ē�.�B9�����΋@7�!T}��ƊCW��Z8�۰�&F��b���\���e/�;���0a�6&$�"]\\ ��(,\H�K2Щ=K4��w%����&�%ʆ�25I.�;��U���#=�VB��°�F�^�ТT�"$�z:�5�:$N�8۝�a.��i�n�C�u��!��5���bJdVݥU%R[���s-���}��\6�	��!�����՟�yR��?_5��r'�"W����=�:İ��򻰨�/[��g��ot3�55R|!����4%u����r�����`sV�>�p'�Oۀ��M�ŵ�!"�8w\1`�<�*������g��W#�^(�k*T������}q�%��w*����*ɸ�[�Vi"J����ݔ�aQ��0Y���ɧ�a�E]��Ο���	I7�:�����ܣ�G�(�[_6Z����X�{j��y˗�g�Z�U��cw�:�1�%VI�G4:�p�
�vy���ĕ
+;��0i�_��Z����6�M�ǒ�
/�<��@;�DݶBM�U_ Z��՚Ҳ]�>�2�amu=!;��1�g����/5'�ͅ��"=�s�k���v*���G�c����9�<��?��O��s�d���m-���}zG�e��02R�R��}�*��_��5q4y5aC���G4��R����e���W̌����������#oF0����~��Y��@�~�P�vrPk�V�q����|
ћCB�~Jh��GO�r��-u�PIԅ��K����ِv�Z<�ʚZ��M��8E��v'^�48�@���JXc�	�<2"d+�c�����ҹ�4�$�{W��z���>}hY��R%��5��~�q�h�Q���k.�y5
��wv�W�g����ɗ�%+]"X����.��MW���R��3vp��t��ދ���T1x5Z�h�n]u>D4�צJ�ۇΎ+*T��\9���}���i����|�|����(^���s#Z�5�]�vэ���ĵT�Q��]���-�JL�/u|q��dKn�bΌ=Ito�j�S/k���E�^Ws�:�)������UEBN<��R��z}�å)�҅��i�7�U��o�opq�q��e��=9�NC���mP��o�󸈫0#׮È�O� �y��+�ֱ�/SF9���c}!ޯMרH�`�բ
9g���(�Ό������K�M�|q��w� Vr��$����8i��ܝ�;��W��!���@#~^���
ǖ_2Y�C�7H��d���uk�B��X��,ת��{�l�K�W)k�mPͧl%��bdi����ң�LPDs/GӪ�t�m���m����XH�v]�&����wS��?7, �=�Y�пw�/��W'°K�J>V��>t���O�	Q	��+��oP��l�Ǘʩ.�f^�(_ݒ��͂۴���9�}	��{�*��1ۧ$�g"���XW����Cj���9*T1a�T�]sv(	g��R�¼h��-\�yA~</GfKO\N�y��O�0����%�cɆ0�A���Z�����G|��4 �Q�W���q�������=y��e�zf�I�\L^jG��\B�Y( /�{�J�w,���	o�'���t��g��j�M��MT���m'g*Qs�6>��"�ǈ�xo��:����sTH�W�l$�{P9w�[�U�Mc6�of�Q�𴮾�Qu������_0c��+�/V�����[�9���l��G��5z*nI4ή���l�<?3��5'��:�n���&�B*��e)�	}�#���Zm��WI^i�a��-�+�o��U.仰�u~�;?ZC���Ĥ��l�
�D��#L`{�s�7Ҫ�b�}(�4^k �l�'[�l��\h��$-Qo2��T6��oe�����+����z�������@X��-�8�]�i�\z��`x�3^#�]Oh�u��Ls�r��X����V�#�w���׈�\]e�H8��QMu�c55dlQ�㫧��)�V�p��2k���X_���xZ�o#n�M�Br%�$�ƭj�V�/���r���N��&�^���mw��*/����M�x�c�cx���������7ڙ���.9������a�k�H�å9/�#p�7&ν�c������h�	o��PO��S!�҇Mn1�B�8W�RH���K>�_�Q�=�׍��Z;#���g%�G��l^)V,����-��yiɳ`N���Bn!G}���15/qCy=&���4�����dM������	�{R�f��Mѫ|���u�t �`���OA�9�wh�P��8.�g��{��h͗���Xʩ~(9��*�u`I�r	YTekd�qA�4Ds����ͬ���	�=�nհ���� 7�{���BU��B�����w|�gA�:��D�l#��t��CIw��ê#����β��Ȋ�e��RM���v�q�gc��c4�3s��^��b���h��n\X�@�5&��F�/�5�����S���ޭ��f������=xr��[���w�i�8��61�����!��6�%'_�kظ9	kT���;���plX8F?Y���9��Ԫ���P���)1{��� ^�YSs�B���2>Y�󎭭�y)-P瑘�m�vcU�c��G�x�����<�q���޺T�5I���Q1N������;����k"q�.#�zzzK"���YQtC7�4ٜsaxm�X��Ƌ�J*��|0Io�F+WԻ���z4_b\�����FH��f��������@1��:��j$Y�.��+�!+���c��ѹ7A��!5,AK_]�\�_1�0!�Zc�q
1X[�#�&�sL�^`Z���)kw�E�W&ʀ�WY��h����,����%����j$�ZV��x�$Er1����.���[#ۄ|�(��p�Y%a��Z��DZ�g,`�q�ڧ��.���^t#�m��'\�4�<�e�
4�<ahZr�
ȝzz�]9�)S,c�(F������H�<�-9hX�aA��#��lT���oe:Z ���9)o��f
X��լ��W9y�^=w!����%�O��G-��8L�����ۡ���-�p_�3HC�� �)5v���9�CV�+ҽ[�������2�S�u�QUz=�x^R�Sc�O�	C��u��~@$�ߕ9���<�?�R�1�	4�d����8x>�Cn�xn��l�xt�7�X�#ӷ���Q�Iŷ�ͨ~mw�ʍ;��ӡe� ����_�8C,���$�4(�V'2�8�hiZ�ϔ��� ����]�Xl���[4j�>��]�hğ�,'Ʒ���3E�+X��ي��uu��k%���T�;*�%��#T6A��NC�߰��kZX��\j���NL0��`r���Ṃ��'�@�d�����\�Z��r�v��%o��s6�g=���K�$,�ñ oБ��cG���[�l�<�#x�y\�(��[��j�YR�b������m�@B֭釋0�z�e�j����ܱ������)�f���c-�<l,Fs$b��7����69)�	�ל�3�7�1�T`��]�.{_h>yQG�2���Y��y��.��쒳��#�|/K�]�cā<����y��
y�~�4i(�@bg7�rYG��N�r�զ�e�<��E^�䜈J�=6��E�o&b���C�[_���l�a+��?+��d���v)�r��k� a9=�Q�
t$"��	y���5�g'�ȘU�ѵ���0.����f�eǎ����o'?C1�.j�o�
T�4켒e�� \����3ɍ��4ߚۯ0�����=�Z~�ϣ�J�0���A�E��Z,�F[�P�AU�؁��*;�P[�Tp�����٭C���)��������Kx�\�ĭ��܋\L��9��ҷ��{�Q\�ّ8��;�Y��<��T+�a�ǛҷP����I5`��������A���v��کk/��o_��Ӹ݃�|T�(ˋ�.�'���ߏO�\#�����{���/!�`��{�a=I���KA��r5]"��.�FJƥ����B~���U��Zv�Z»�\�8w ���U���9<h���c��ނ�ԓlmF����	Une�������W�@!�kڂ_h ي�ra���03/��w�����{��U� D��rg9�D�~2x%��������@<��T.�g�%�/L����4�`��S_-��^.T���ު �9b�8��� �����tՙ�z|�A��*r�4u�7g�Z�36�7Ns�]f/KK�X����2i�o �xy�d��0[���Q�����L$Y�JG+i��EP��9t=���r�k,޻�2'�9݋9�W]ϧ�`��F�e�/�:a��z�a��Y��w��5#��6���O��X|6��=���θ
�@��Rt�W6р ��Pէ���٘-f�����bV��Ǐ��ܤ��
�ζȖh��I%��#����*�PY��6����X$%�{��,����R��C��`zV�G�b�:�1X}۞�~5�4)XSs�]~� �|��k6D��,��R�Hҡ΄Zua�@�D��amHUE�9��?��A:�*�hQF����^�a�����@X��_f�z7a�k����ـ����d��D �#�h+��0;+y�tLP��֜��������0���.�w����m�m��}@�>���ʒ�wu�Z1����.�[�W(�l<���?39��R�j�{���Jl�����m��׉�%BCbZ�AM����D��bS�*�u�z�V�q�5MBoRԕ�,{i}ix���İ���~��'┋Ͼ��<���k }�j�Y��WGA7�݋mN��?�M�B���[Z5!�4��^���9���`ԣt3������0�z���a@��P\��bsG�����ʂ�k��H��<٢����`xu���|�Q�R�՞Ae<=3R�&�l�G���}Z�j�M	��d�@�"��Ճ�CE��#��4ݮYH�K�T��zh�[�J����(�p���7R����*��m� ��17M�Z�H�2am�O�����1bq�$mc:G�Ve�sd��."L�G$UWc�5��4��!lY�Ӆx|)� )-�<|��ǝ3"Q���C��[��Lu�B7�6��a5��Nꌊ��J���a�4�3�uQ��bQ�yM�e�����f�95u+�x�����h[Ȝ��㒪��5ԵӶ[�Z'������L� 4)j�w��T�J`������1�2£��uO��Uq�-T���Пcgq�;LR^FA]P�ܝ�Ea���[7��_L̟\hԲ?_m��c��EGPO��)�h/�*?�GF=��6 �ҡ��ߪg�y''?��]6��ز��73���*"�����1+_O�(���^�i逭���/�h-)7�(+�����+;PR�.���Ц�����7m�^~���q�7y�j��X��G��!����?��M��vJ�4���wu4��C�j��2� ��>t��7Q^@Yʻ�ӡi|��v;��>J��u�OQ3��5sV�Z [��j���P(����
br��ۮ_`��vKX�C.�Dc�gC@r$�IK���܊��D i�ޏl��>�@u��"i�/`�k�qg�d2��n�G�j�5�(vv����C,P����Q�@�5��	F�7�k��Ҩ�v�A�?X�vg���/�U� -_Mwܑ�7��op�����@��u��	M�.���<�ܫ���5�)���F�NL	 	�(�F˂�2�q�G�W�4����0F'48���H�`5��V��YTl��[���Tax!Ǥ�)�����R��(���?RQ`�>�q�`�a纼��]��.�՚�p

��J����l�����+��/\�Ҿ����L��Wy��H��Z�R�������J��ƨ������v�+�[8U�V�Q��)/!=�5ש��N��;ŧ���zm.�L�oB�Ӊ+�f�����A�l�,��3�i��ã#��WR�>I�3 ���9�$�h͈��O��j��VZhC����^~U���U����ZH�R�3曄'V:�iW��}&�Y��Y�^,�,��ʓw��
l�L����G,�l�	�1bN��&X���kX.�?$x�@b�%P%]�TO1�����P�ˢM�k!���[�^|�;<�I�h�>p��͛�;�U�RKv6�ޗMO��yj���%�K�.cP��k���
���X��]u@P%���c��`�P�%^ JH_�N/�f%�i�q��Q��,O�q������+Xь7�/}��3A���iɕGF�}F����S��u��rer�$y05E���kt�'MF0���l�F�N�v�p5�l���.0��:֬�S�霐�ˍbz[��bH�E|�^	�c]�,P�3����6:��R�ԟ&=��ZF�5UC<�֯_��6�Ar>}u�-��1Jڇ|�㿖�k�Ԣ��ÏT[}��&����4�&��yR�;}ݨ��*�Z[�e�!<i�+P�P��^*Zhw�.����[�f�M�識�1A��r���O���T�r8Y}�ՏP
k`�@.��q��z�U��(f�'�/y��<�_���N E @i����J�אռ����K��H0�m��x�����5#t6�L�
V�淐����8Uc
�8/�	X�.1��h�%4�Eh���v=����g��2�6�Թ�q��=L��j�FOC��4��N�Gծ@I@�@`@]ZI�@g�ݾ�.�R�F!շ��V�=!�#@�^tC�����ٍM:����By��$�O��(4h�n�"F�M��N�M���lm�[E��z�:��%��}Y/��ش���9���R�H���gh�!�t�w��8�D�fc�w�q�hrv}���8�Tt�q��>��V�S�>S+�k�	�Mvx�7֥`�Ɉቘ������Q��U(�!�I6[��]��c5��_�ʷj��j��+-�ǫ��9�.>�幒��s�0�YB�JU/�K<�ڄ^{{����(���Z���4����P�M��\�`6�OU�R#�.�+����©�c�%WS����,K	�m�C���L��U+*	4�O�Z?�|�8��_w�
��+��\aD�I	A��������ܒ��|u�E~?-�Z�Bu�6�A\������H �/#s �W�ďjjO�x�vO��k��7���4�	���C��ayD�6���Y�d�����'Y9���q'p��z��B�i~���S�g�33�x�T��%���{'�!j� �O
��9�4�l�B���Q��V�w0�`���Y��eM��٨g����Қ�Q��'������^g����Åѣj��K�=��j�#HS�����"�!�+�;�N�`W�U���Ĉ��D'���-�r	@�ԓD��gG�B�\yWԳ�t\����s��~cE���'*3!ސ��4�pѤG1�8u�^���P���!��e�e�k�a�9���þ��l�~.Б��zFZ��T]i��+��τ�|�
�R�I2alY�_�'��?$1 dI�92n|VVǨ��-W�L�p�TT�)<��xT���]�bƆ.�B�JHN)We���{�%򬩥�i>^П�E�a_�Ɖ,�Bi`%��ƨ��U^}S���oT_�{��7�J���-Z3��{}�CYAt~!|��Ja��`y�`�R`�S��]3s�$�(��֯_>�6
!Tױ5aa��1�4ػ'g� �t�_̛�=�����v�u����v����gl@����1��*����ꗆ�M��0�[-�lxA;\���`ݼ����1�|p:H�]5��y���yŚ`��GkLô�a���O��m�k����13JқC�Z0G��RG��e��������D%Y� �77���gxAmWk�!���/����g�s�b��8W�|FY��7�%b���
����X%u��>,�֍�_&:�7R$��zt񵒊
g|�u�=䒾/=G���������Wm	��=�ԾR���RB/%;�d$�r��s��JO,���澄��ڥ������;F�`v�������/t�j��+�a����{���_\������_�����g������V�Ż�7PK   ���XWC��)�  � /   images/093f54e3-331f-4155-80d0-fca9fbcaa25c.png��	8���?>ҡ�)�T�9�TBC�,5��A�(Kd��/�q��2r�fP1ɞ�0�Q�
���=�k�}��~�z���������{����y��{�_���ǣkښ<?���\�����.��~r��>9��"�؉���]���u���K7�0ؑw�v7����0�='k��-�;0��v��h�[�wN;��ď�?��
����O�h�O� ݯ{~bz9a�.n���(��@�n�OoF�������_��v,ȋp�qW,��!��U�Է��N_�W��+��ޫ�}���.}�s�����}2lTSr��i�� C�s���sJJ��i%������鮋��?�������� T�źȜǾ�'w��A�t�+��OhEz8Ϥ�/e�>���e�%���%O��'�3W�L�����TV^&�o^����{��b0���.+Ű	�~�8�O�m���z�K��n��矌�t��d�D��`���JJJ�a��8�]\o7��N���;�Y��Kxrt�
Q����G��jm$M�KBS�='{�VVX+���i6=�˯�hT��_�1g���a��p�ݥ���6zC�*��4?,V����U�\p�{�3xc�w
C���\�"��	Z6�{��O$�O�(����Wj%�X����K���}�u�=���'�5�^%U_��~��!a�@G����1���̦a�w��W���4�8�$,䄞/���v�G�����^�-^CY�	�S�	�n���!T�17�!~,){$'L#Y'I�c�*1��9H	���|$��~��P�M�P�?%ͬLZ����{�OY�'L�oUۿH�H��������e%���OƯ���CkBW���Ou����Ƥ�n=`���C�\������Ŕ����ORŖ� ���۟��(����򣂒WP0;��e�*m>���G]�
�i�jl喨4eX���[\Hk��������6��ņ�\�B�m;�=��U�C�89ݻW���sv�~7%�f�J������n�2�oQ����u���^ۗ��% �5��£9�Z��;��� �1����p�`�g��7�Zt��nf��J/���DvE�.�5�b�`=ۥ��"֛�����K��ͫ��C��zCq'�sN�z�N�����j&ӟ�Fs�/��!�;�p�ԓ��8�L�aOǆ�{�����BT�}��dPTbߘ{1�K� ]���`��8�6JqSV�K�O���0�`u'��oB-¼�E��a��+��G���s�.��/�2��|cB��6]�`�2{��TW��wAR>ڦ�ªIϕ�s��}�z+/��Ra@�;�b�.NӍ�;n�`y�O�X���V-M����������D8`y��<�D�Z�5����`ҵ[���X8>�Q�+�Y�m�L�Cp5~"�i!����a�
���	�MO�����B�"��2�T7����\A�I�o�}8�àq�`_�K��w�.N��<�_��r+���>�m�0!��	�?���c]dkjd�9�f};OA���HGX��[[�klHR���B�I��N�-%=]�$X�v"ɑ4n�<���v�{Ы����1�����m��(�_?�'t_'s��n7�Z$qR-g�}�����
�3�U�	�ۉ�Bk��c�4Ƕa��?��d'L�_�� L'@\���P�>���u�y�f�O��1;arQ�	$|I�KՎ��^nKɳ�4X�,D�|��"93��"���$�7Y��y�������@�N�K�d�ct���}u-�D��g�w35_��e� �2ty���dM��E�Uಷ�'�;6>���X/�I��>�ѱ�*&��7_�~7$c[F�O-n"Y�'������N������-��C�*6g�uv�����'z
	��r�/@B����p�\j>l{� X��P���z8�&7/o_qq1��w�7~Gg� �5��O�|��Ijs$����md��41��=�Y���E"��ll�]��wӵ��x�aΗ�����b���w�{q��lO��5ޣL��3ZVZ*���L��6C2�\0��`�}�^,��J�t��B)��x�K��x������$zU׏׌<`ۋ��s�.���]�J��ˁ���#�9�!@'��q6���$�����/%e ��EM���ˤ�(r�1��zI"���� zZ�	�����߾=JM�>����WW�e��Y���9m[9L�(�������[��K���G---����f9�1{RYQ��&c�.E}9�]�Q���{K�r0?��%2�%�:^3�YO����?��dH�UND�k�@ �lz����S�9��Fp4�����h�]�|/�5�_DJT��'A�����^AW�H������ b^��z�����z��efeU��Z�D"��e�wI�o���Һ����%!��k�K��n�^������rs;k����W�+���Ȉʷ��o���MI���Z�]��󘻕���w�C������FF�@s�F�j��[�,�HZO+�qm�n���@_�w�{����f���w�_��6r^�@�I>pC*�ӱ���q;۞=�)�@e�A1�E#I���+k^.uK���'jM?f9� 8�� S�@�T��.��w�=��U]dnI�p���{��%���kS_���S'(,�Q	f��.�����f�kn|���Q�+#��
 ����g�T/�����Y�y:a�x�[�%���*����f�4UQ@!/�2��p����W'Xk����u��ӧ��e���[��S��7��c}:[w��1��rv6�b𾿫�a�g O^k8��<���f�\^c\�s0���Uv��w�
ܲp��V^w�� ��;��?ݨ���MC� �M:�M� C��},\K��RZ�B�&� xVZPp���X�{��E͎�Ύ���S~�=�y�tWj@�XV ���<G ���ؓ1�;Zv���5���Ά�V��l��&Z�	Jh�^��kd����o������������{珰���6�)���i�,w�&o�@�X$Pڡ�� �4���Fe�)<�8��O�!*7141	u/6U\�� +܉i.��0��O� ƺ�:w���f?^7�^,sp�f��t��lhf������8U /���@����l�T�	�5��it$�ޘ��%�O)>������Y{�h���t�����	�m�ja)P<͇]����(wY�o-yꔧ�Z���x�[�'���<��G(�mm��	��X�����Rp�[`)}�ROG�H��F�E�8�3�	]��}��m�L�Z��k}�ES]�w�hA�r�����C��ќ����.�&��-uC����|7˴{a֨��fvXq����Ps���<{�#S�Z@�S�d2����U�%V��ә������q��������^}Avֻ�s��j��A� ���f��U�(V_�N��j���3E:�SO(7�|0��5w���P\ؿ.,<�<g���� ��Fe)�X+H$���4����F_YLb2���D1�_ל��.
u�ԩH���gv/V�O*����w���AS'��EA����K�W�"i�Ts��_Zzz �XPP�'f�V�u���7��:EvQ��~��}]i�Z���{��oG�+��C�3�p��HF?v����;<=�Ez�����&[���j�����$]�A~~<N���ie."��Je���]m�=ɧ<���B��p[��k(���Z�g�_ou��Cj��Z�7�]��:�/EEhV�Y-6��L �W�u_�X��M���y��J��z�k��/-d�!B��������ۤ�3�6hBU��]��4�,��� ��%���^�B	���������6�F���ă{��lp�őhF��Øq��~�,�G	�k9-WvĢ��p�@SμL]��.�bU�T�99b���}8�u�HrDq����\��j*bcku�M#�� V��Rh ��qprR�z�"��ž�AQ��ĵj8�}}�EW�#���}l�<&�8�Q���xr�wR��`��Mӫ�
�A�M��(ƭ���M���o�������)+۞$�ƶ��J�%%E�]}SR�;j���oԦQx�])== &8�����)�J���u�rY�o	���Wy{��_�r ��Y��=�6�WC��U��<�f�i"% �k��3r�"�zC�����gC!�,�J��b�~�����������n�	�6tBHB}��z�����d;����8GRdg�w�c@��
��l�����0YeNl{JJJtqեӭ��d����(�ȧ�����tl�3�l��vd�gS��J��I3����?ͱ���6m�c
^S��IV=T���ODy��t_s�V
	�]���+�}!h͟;Iv�f�B]Gը} i���4">�)tf����<4��:��J�'e��-�([.��z��.r�)��M�o �0d����wHGܚ�/f��?�T������K���k�=�����o ���>D������C�5a�]���+y��_�������9�f��*�;ǃqX�U�^MO�p��L_�6�p��͆7S��> H���j�8}�N� �V�5���ւZ'��QH�������9����Lv{�M5���;�]:m��{X�yx6�
�U���ꦭD�X��l �@�T�D�)�]��<*la�PWo���ux�j��rF��!�Ne^p����O�̸�t����_�YC	R4���&���JJx�Y�.E�ɣ��S���p�j�T4�J���қ����g��.�Q�'���E�'�Ν;WF�삭Q�f�j���1�6���ک�<�éQ� �e$��ݟ	Z�Ys3��@%�-bz:T�)^�/��~q��SfK%�/��^6�ʯ�$�DY��� �O�5쳳�SF^Wm�+$Q��\n�$ �k��#؞������,��I�#����@+p�J�Ȭ�>����"̎'�~�����o�ċ����GX;]�z�@�~���&_֟˝F�49��Tzϒ�V�����Y��s�3�g��`,�H���k��yl�=���9>�745M����j��Ry��w�TB�M��	~�[� ;��`�h<Zg��~�v/wu�4����6Sz���J�$�ZҕђH]�t	�訥#P�>]�?K�����V�Q�;-���RampX�Ř_ާ<Q�hߤr���R��t�lΣ��D�Pܪ�=劲�|�������e�]��cl��֯�R`�,}�6]���.��Wf��\+x�+��W���s�Sk��q,���Xwi�Fc���}Y���l(��+��O$.i2P9ި��҉0r���#�h���ȁ��co�M�͡O�0)�J�[��� �������𝮟���S0x��1�a�tB9Ɛ�`�G B�KT��Z�� ����d�|I�u��]jDؿ���*@���v;�i�U�2<T�}�rjk�e��i��������Q�+Aw�&�e��=|2;�����R\Z]�:�$��@�%�1�z۸YV�(P����Ŋ��],�|M�G"*��q�j��r�J��,y�k��䐐?�#������������&Y�]^U���3�8^DO,y�w��\����>V�<߱���(�@�ƠQI�k�,�س,//����,?%��1��˫h�g����Է�S�Q:b���n�s�{�wͼ\h|�"���I��)�i��+D츷��� w�Ә�i���kÈu��u`�����$���v���-T��T,��UE�K�X�Q���g�P�A�fؙw��a2@_��5��8�'�fyՅ� �"����ay]>�H��'���$��[��
&�Z��}��*!Hu!�s�x�h(��ݾ��. h�P�s�*?��_�u��Nm�ݝ�~�C�V����������W5S���7�x�L��h��TE�|�A�����A�#���'��ݓ4[6�Uno�vB09;���L����;��q����d�I�H^�77��7o�G�z����O~Lf]g��&+�k%}pM|$��KM�'c�Ck��Z)G��B��Nii�E��ih~X��|�~v�l�r�M�����J�p�sM����bta��I*���f�����\W��,�c+$M���g���Lk���6;Zq��ɓ�c��m'&&X��o��[�VL.��dc�)-���%���w<���n:���R��l��H�cW��)�M=5��KA8�{��Lj��r���s���$�}a�֜_�  �S�O��w��>�ɂ��B��������5R�Ua0B��[�2���Qq�9�#�o߾eZBlL��o����/ �����������X����gO�?�7���_6����j����H	�xr�M¹�-g����3�ƿ1(ZӨ��i�#�X��IYQi��(�@+h�X~����pG��E��֚�(TU[�ԂH�}���S�F^��<?k�PEU"=[+~�C#,�\����RqQ�M�\�O�0�
){Z�5_������֞���V�i��mvv��	��bd^��I�ø{n�x�|��333:P�����A�p����x(ӎ�����AqmN;UO��	j?p���|`�g����� 5aW����'?p��%o�
MB��ϣ}�`FisؾȚ�7����nM�brA�
�	���/t�2¼}��Y�0a}$cIS�o��t��R�A�(�6���:��� �<J;�d�X�bB�xZ�ܜ�_�OhP���=�oI$-�p1���-��'� �"�(�U�	]����^��9hbs����ؐԶb��:%�ؖ܅?���A�TS"�n�i�'
�P76+=�-GRr��fjs�U$�~0�&��X ��KӻZ�>h �q@�=������J�λ:�A	����
b�<� ���ݹ�_[|�E�jf�)I>��� ���U�h	$?qq������\$�[�W�3!�d�&<f����Ļ!������~qm ��6|���TLX)���<��Ьw�?�-�x� �1 ��!_���C�p�r�~�M})�y8�7� ���;;;i7����h���(TPAHK?��꿇+�U:�|R�(��
>8?]'˞Kwu�12�~��Bo�m�C�O`i�;��@��:نJ�V���#1�!����>��2wfD��t���^��s���0"�Wh���[�m��W���-��!�`��gc����ŝB! ��84s�*��IQ��@��8Ȝ�995iz�� ج��\ޒ1��o``u���o�><���[�hȽ�����M�v�@Un+|��Ǟe��� l5�ѱ1���k���aY��T78VFy�����/n��R"�k߹s�#Z4�4�R���c[^t�BF�wS|�#I�n��Ѻ�)
u���T'S�6����w�0� �����/��h�>nAd������?mP�}���M���㝅�@F��&���{{���e	���Yb�����A96�	��='kYq߶נ�2��7��(|]�_��J5	�Om�����r�;G�����fF�6�]��+֘��}�H`����у������O��(t�?���̗���vh�
��2��/��
Ƚ���p�߫�NG਴CU ���{"��`������z��7\&;{(�t�u��V���D��+�n��SRI��R����n��}��V�翐�����2gA���r_:p��(� h���A�@�5T��.�4Y�St_��k�ׯ�����`	���F�s=S�a@_���ͧl�����9�k�f
�{2��Z)pڄ�"�<�ޅ>����% A�
��i�t��rmSu���QI8c0TT���w�}g�w�燼*�
��]MG�A�(�q�F��IԂv�<'��y�%l5���l���b�V_�P'�K&��!r�^��%�}�i�}�=%2���Ջ]{_dgqx�>/���TF��=���+��z��h�s�n���w
��B���u�:dt�P��x:����ms9�k!�t��Y��n���c�p��ۭ���T�is�-���R���w�@mԶ=�_V\�x#�[�-����������`�ݸg����@�b˵- a���}1v�bon[�]��_���&, �b�a�7�I �Љ��	� ����
����䓟�1j A7Q�Y���F���Q�(рN����goG//L�a��� �,�g���:8�uX��7����{9x[�?<�z�>�/~�s<�?��m���Y]�5�/L��<�ǲ��o��oT���u��������޶G�8K�6�.�f�l�W���t��Z�~���~�F�����ȝj!�FQVgdo�S�(��(���y����e�D}z�CдI��Kg�˶�I��k���/�������ہ���@���o��ÓǠ�`y���
����}y-nVm[qLbM�����A&)�9����I�������.4�՝��WĦD�BzDm���5�֗�.�k�����z�e�� Ɲ튌)(2����5�#=@���S���hZ0C�O2VO#�n���K;�T����\�r�޼��w�rq���Ѭ��e�D[�+�ڶ����qO"M�-<�}���L���]��ҷٗ�SH��^��ČG�2�	�+[��H���7���2��;���S�mn���4�͛�O �a����.<���8�~�g����gB���	�׹�N������oR����,L����O��Z�4{��/�%on���3��E��Yږ������:�z� xݼc�Ti���%���JܰR g̚@"=�o0IB�b6l�켖A� �8�z�#L<ՈY�:ѹc�aa��@\˨�V�{m���n#V��x��>���<K��au�h����d�gu�;u����8߆y^�"��@�`���T�1;wI�/Ok���B�Dܐ�����_F�z�!M.��u��K���r�%��OV�Ն�*���	^��~�sbp��&Ӊ�i�B^Se�}�q ������[���81�ǘ�DM�"�D�w��Sp���G��D��D�����)��4�T�����::2z��� �1/yN��1i���3�1��!�!�?"񗈤��}8o�5����5(1H�(��f�����K�:���r�W%��TWDۋG�(��^g��º95�dro�N�Ж
�
��D����!_语z�X~�F�p"�^�h4;z"�&52I��������F#%[ \��Ng&uY�u	3��UR������j�Cʴ����kJ���5�Zn�W���O��T\w�B~s[��r��h�&l���U0�ъ���������u=����(�W����FVrp���o��M�f�-��{_�:/�K*	��	׺�l��&C灧�������}�����*���j*�uը��ΟF��1�_0li������O��2B���U�e�St|��_�m�+��;/�N���L�X0���U{�ét�V�Kx��,|��/Q���W������NiV���)��;�TV$&X�q_gʗ��Hʝ�~���{68/'�^��������RC~���p�LnE�����bt�%���qF*Ӎ��Z�EK'�7�\<-ֻ@��ef(vu��ZYmyB�'_���Ǵ�3C�n�S�O��J�H�g�B4����,�����n��ު҉���[� �=2�&�mU��}�����_%�)��	��U�;����3�qY��d�OUg*�?:o�\S��w*9�Zx~ �q3������%��r�if�W�x��*o���R��	!���)7�/�R����Z�vJ�az��a��V���H��A�\�~��Y��vإ!<ĳ_wΡN%f�W2�>�2����P8���`��o0�'a��_3f�P�h:W�6�	�(�k�2v@5�?�4��pd�!���X�����VB�̡���&U��Eդ�(2S�?�McPi�U�2����5;|���&�-�P�њ����+�����4E\������//	o�+�Ӕ7-xj ��_B�*��f�/�;�yd"y�S���Ā������1�q�ܚ<<��Z]ɧJNm��ޯG��9�1 �I��i���U����y+���Y�j�;����307MU����#�(юYK�����vO�h�x�S!񥘘��~��WGK����>
��$���m%�JB�҅x9��f�g�%�iz���8��-���b���fi�����u˯'Ȇ�/7=�ߤG��i��؊I���6��ϴ]jiӸ�s�_�ߌ�Q+��<3���8sO��ȧ�ZR�7\���q�c��*q���sZ�����G�_O!����5~�z�Q;)w8y��Hd��O�o� ��9�S��&�v�`^�� ���q���	�#�m淪��[�>�4ɼ�(�$PwA���� &�<H���rƌK���$� ��.zJ�C�G�m�߿/�3S&�o����^Xs�>�t�k#�}V/�\n5����X�蛺4��)���+�:�6���������¢':7����蝈W&������H��ԒK�E��R������ϻ�8��\W_�;Ж?�������;��[�B�ԩ�)�Z���R#_�g(��dgg����S·"�O�i��vE���o�����!1�1 ����k�_#����{)w��-!W^J� \�#��#�EEýK��i�=��/]���xxh������i����[`糼�^�o�0�LMIe��Q���G"��ej�I�:��j�$�]ۓ���QQ9~\�i���8,6q����GDD�p@�Ѯ�Vz���сJ�c't�U�ȫ�Ȋ���ݽ�|�U�ik�x�u��]XEj����&�ʡ!���P5���p��+R���ے��(�e�Z4�@c��.���D~e�q�#պ��N��>!���n-�șH��<:�C�rr��� Ä���_�E��'�L22��<�>>>Z�� �A�a�X~�b�S~J��z�~�E��L��-��&V{�Aȧ&����Ԅ�W�����.���_��4d���zx�ė�i�ɬE$�D�듹yմ��x�z"惤
�4 =dm'Iihjj�^��L"���T���nH���{%a�T`9�O�R��7Z^u=�U�+db��C
����A��6NJ��=����)4,,J;�}�[yn�۾���p��U%^�Hq��CPV������OR$��mR����o��`���JC��-�H�u�B+F��Ç6��ꁷ=x� �,u@�L������ᝃ%�vmc����c���O%8t���������^?�����کS��[>
y�F��25���hW�ҁ�&
�^��lfC@Ǐ���W��;�|H��ڝ1Q|V?ʳ�q����9^899���Q�U��}�����2��3���v�^~(����&���j���v��ỒWJ�l���)�cv��L�>���H(.X}$w8�������`"$�B��#w@(��k>�cZw-��"k�����bm�%h]�E��)����ۿ�ل+�У��ī��-4����5I�Y��tx�+^'ܔԜ�4S%4�5
����l���U-i| �L�����ӻ��[�|0�	���c����\v���ml������3N�_��Tg�H�UY=����4E*��������i{.^FZzom�dHYY켃k�<��v*�~F8m�W�9�4���1��o%9AϿ/��z�Ds8g��,<���z���4�A*�v�!P��}A�!2�Ǥ�`)s>�7�����W/N�ʥ�:��`�5Oԇ��ntGC������^����T�������C�����R/�@�o&��k�B��7
��D�7��[�tᲄ�)䬧�|�����7^5���Q��L�ʕ+�==��TL>0Og��+5�6B����̺���3��.M�ូk��ϯe	?��9O�o�f�7��j�MҎI��sc!��ă�+���/�<9�~�5�+y�ٝO��3�[;ᮊ٘�j6��~�o����W-ws-��E� v?�[e�|���B~:�~8,��*mM2���j��Cg�(\��H?i�C�v\�+
�#���xEnX /@���-����W]Ԧ������ˊg4����?đ]��=�{+7:��z/�Fr��3�>��@m�����ſ��E�eu�9^4��l���V'��s,[i@ἆ��@������"�B��?<||��fR	2��+[���Ow �pRj��w0_�m+�vu�-+�i�2W������ye�z��g��Ď�I��KO~���a��WJ�yp��Ԩo�Y1��`��%2��Ǿߴs�=�>(�"�	���o��ci ށ;!m�.�J��e1�oAߪh��0������a)�.�}���I|`�(X��8��EO���&�0zéVׄs����gϞ�
>Ua>�g���;���VU�����M��BӃ�!D���7wj-�����9�K[Թ;�U^�	+� _�q�X�AX���\Y�mydW���o<ԏ�>�}�z�jk����-�!�6
5$�ғ�T�1�8����"��pE��Ґ�`��eW�W����ŋ]*�5Ր��iqB�T�2��=���f��iiJ���z����&#���/���[��t�8��M��h���#4����Bv1�py�85�����j�Qe�ѹ���t��FE6q��^%S#����56==���S!��M]ş�Պ)ȝ0�k�B�Wͥi��2�u�`J�篢���w�J0S0�Ƙ8]�gnT"a2vy���>�q�{u��f� 0�|Z�ݠ�k���0�R]أå����������N�i�c] �02�	o�./���q�i���ʒa��4悙J
�Sh{�b�l�Tr�5�����dIř�W]�����bk�@i��4_͵��+|�{_�bֿ�ߑ� ��jqj��[Q�K+s��AE�M,�E���Gj#\<����0���dM��ORV�bJndE[U�����<z�h�A�/@&�~B�[Va�X�>�n�mE	�����:w� ����d����:.��C�K�:t���K0�����3k*I������Q$��󱀹<���V���R٥sm_)Xl<���QU��^Ԏ�� R^�,g�[���9���,�J�YU#�b���I�dA�;k؜UDh���F����<3�<��6�;�G���n��$`F11�**��d9�%랼#��X4���f�;��86��4�IE�A�to�����k��"�4�	�E#X&S �T��鈂�j�����j��h���¹6����� ��	�B�.O�-�DpܕY淼�/�����߅�' o���h!�A�|������O����m�h����v���1�l�I�72�m�ւr��� ���A�4q�vg���/e��?@�k,�ȵӻ�����A���3Q�w�Ų��	A����3�{yL�5zE�������rT�����/Y�}>��fZ	����\bW��6ߦ��ʷݎ&˙({Ǒ�H)�>�'@|6����a��E���Ϲ�X|�AW�m`n[���;��Ż̶��|��S�Ar;�Sr�
coǼo����щ��]X����og)ͦ-�8a��O
҈ޫ��g�����|eN�K��%��ǽsg��P3uB�����V'H3uqg��&.� S������P�b��%�M(�P�#R:��m�"��j�I�<WU���d�WWpŃ�-���ϗ��r�\ANU�Gw'M֦����}�c�O w1+A�m{��ܨ�dNz��D��D;j�|�?�����$/:��4�d���������QN�ϴ���Dp�FJL̆mJ��׃~�����5�ة�RN���
����A��j�F���A�e�epϘ5�H{!����]�����"�&z!��#�1�/��ѲL����k}�F����KJ��'�K�c.,�\ ��'X��>@|�Jy-P����q��BG?���(\�j+o)��,�㥩G�LL���qI���1���t�9B�%�Js55c���V�<K�R��H�"o��E��B��zsZG �7r=P��~Y5d�eU�Ĩ���G!�i��P�J9;�7-^.	K�Vݲ���g���[=A+v����|ױ�A�7�o
K<iw����:'''@����4+%����U�h�
�n�T�?O:)��U�-�}XT�Ջ���4i�_�}�k�$M���2J���i~�KX��Ț��$Kޯ�$�H��t��+[�"��O���r�xaԾ�����M� �h�H�'�,KF}�Ň�|��kj��+F�í\oV��+���g��8��(W[9.w�^�5�Dݝ|�ar�y�}M���Fg�E��C��ے�S��.�����ch٬dNNN~@h"{�ы�؃!���e%��_++}��$`���i�J&��t���.�4���_X����vZNR�>y1�iL�!T$^w�'��S���\	u��ŉ�!ϘZtG�4b����Ȉ9�;Ӥ���Ғ�J�w� ed�y���a��9=zd2���ZZ�6KԠ�H�{#�I���T?98.)D�����J�s��sj�����{��.Ȋ�W*�.w,����/���A����B���͜Mjƃx�*M�F�4�.���냺vtl�@�'IY�B��
fw�u�neC�X�:V��wv1���쵻������G9��W=A�M��q��-F�N4��������Y�ң��VSID�)@v��}�+x��F�}��=Jfe�1�.�3��,�^�tu��#��w~R`�W�WAAA����Š�ڬ�� �R�vQ�]	T����6K�Ɉ�-T�$/��<�]�Z�ዬn��IY�?2�����!B��e����<��RDc}��0�)���볁	����>͔H�z����݈׋u������n�(T:q��C4�uh�:�CʩM�u���\��.����g��"��U�!(�����Vۣ��0u�L��Or��Ԡ����~(��E�]��>?�i_��r�k�w_����(F�.6�t����'��(k�X|�o��꣹��A/d1��b��qMh�԰�ǡ�
�\��#N_�?չCR� �E~s�2U��"wl���E�+�_��Nl{�����s(��<:���2W��l����<�rW)�8���D+V��*����Y�� ����v;!1:�0a}�؀�X�|��U{��n��k�j��XYN�p�oO�.��EZ����]�B�ռ���uv��&�3d�5��+�����\��{��*�WEn?V���d��k�8x/U��@r���>Wo��@�ӊ=!"�ǫ���o�"/��(ned���7.766�&5]6�d~X����Y�ߗ/���m���c"9o��d��"�1(�A4�= 2� "E~m����ņ2��AYM�OX!�u����Hƹ��e�Ӈ��V�q��7�1�m��W�hD�+��B�=tas	����Z+��l\D>��-#�=o���*�0jݏ�W���_�]nr#��RQbce�c���Y ���\�:�eu�ۄ���?$ٹ��?��w�Q�0K^�L,&�e���%�n&�7�&����f|X|/��I�����1�sf�x�?�v�Ӈ�m	�e����~���@�/���$���Cm�6�G3��Q5Z�n��� c���������F��V)�Ŏ��Ģ�����9��bE"���k�j&�w��cO�K�1��W�'�N�}HSUw��I��|�%z"ᬱ���_:���u$U�Å;�(V�~�Nh;l�X��Ԑ��P�F�YxΉ���S��.~��*��	Ct�8�2��s�X.j��:�^��2E:aO���R����a�T��Lw'|�"�l�i���gɵ�x��'ѣ�6��FW͜qd�F�i��������x"2�5+Wh�u���Be����I�t����9�VkjMt'��V�`�(�@ݻ��#D�:�C	�4�
�:���=4�N$T�>;�;	O�����)0�>r�����+B�!�ETz�gS5����)/$P	��&��d�;.?�;�B�� �^�_˲anL��)R{�[,�+5��g�..
wSn}w5F����9�:���u�q�%��SV��Yw� �,b1P0���r%7�&�I��5F�uZ\W�����6u���3���4+�76��,�p��O�C�H�x�V��[�>0?sz�Ze8� S�l�jh�v�@"U�Xw�����S�Q����g{a=/�}���É��R���=Δ�/\�g>�`�s����Y �_���.���氂>L�ý�r|~O������d����Uo���]�+E`��E��@oյ��gJ�@��F��g��!�BWz��L��m:�6�~�I���
q�H�.]���y�ń��v���N�����y�� ���/L�0}`� qD%z��,�r|RG�\pĖ7���yN��L��˴J�T�ӝ���)�o^S_F�j6�����$�OƎ�B�~$��E����a2";��T˓�,�-��I�Gx�b���i��1U[�d@~*��Ŷ�wM��gU"�o
����T%�O���F$���	������y����'���e�|
^�߱@������k0/x#<�g�}�O;!����3���e�0r�I-"���/��Ί�3�>M�֌��>��r�,�;E���O�^� J��!�m�mï��Ὧi���䊹���W����RԽ�r���/�%��^�d���v���K4�w�n���Ga�wX��dH,Tt=u��O-_Uץ�����5v�l�.ߐ��X�u#{UF�Y��1t��'럯���:�T��ax6Y����!��Q~�`�	�1�٣>�m�Ŝ���j{;>�
Ψ(�;g�Q���t��D�^"n�2�V�}��1 ��Y��VU��a�yNJ��(ލ7��V���5`o�����_Ƚ��Ӻ Ü�rk�0f���Mp�ծ��U��2 ���jK�+?|HIo�21�G`� �5��}�Ŀ(J~1��I�m����V��j7g��rY�|2�M�s4E/����#�/���8&�4�h�|�xV	;0<�e��4t^H#����Ǥ�)zƫ�ٹ'Rˎ��o��!D�T�����_y��S��&^ܶ#д�%�꛻��7;^�`�V�z0Vy9^�6�uou�rj�]"�(�8�V�V؇�1��������}!�s2l$�,���ů�x���}%q%�zl���*�qg�>vr&�i��[��5���_|ഉ1��U��&��ZϠ��� :2U_?��� -���	N�{���ݯ>��?���'��~Ǫ��'���A����E+S�ޑ��#�+�)0{yJ�n��%z����8�����x@�p+��ƿ˹\����8p쎎6��^4�F'�w�cO9Į^�cr�%J����^�~��vz.{:��f��9�St�J
���#Le�G��H�6z=n1��o�`W��+o�g��"�<���F�[��;:?U�� �˒�|��SRxv�y�Ԭl\R�AJj���nN���(rPG`ަ4��p�ʤ0h0��px�6��§�`r�u�����mv�N=����O~�)r���e,����.a�����O�/���W����m�@��3K�W]-١»�$��ړ��$r�nm��B<��k���'f�إ&���jx`&�_�R	݅ ��٬`�p�C?��=T�=*��$��.Fk�"��#
tJso�?9�j�y~\��YX>mR�i(�ab�A��� �~�����C��9,\�t�)���>+bƺ�F0R��$���+q �����Ҡ�!
��6U��i���vI��Cv,L�RlU�EK���X�e�o_A�~�>6�ŏH �Ib(qTrI�ɶ�FX��IR�\�u�|�x�ͥɁj�1�-�a����h:��������,k��AP!TwUP�"]QP@Z��J��KG�zD� A:�C�	=@(�|��Ͻ�����������9s�甙9S҄�{�|e�A %v��=3'<�9U�ԒN|ќ�nM��XbہK�ڃ��,�ӑ
�w<7�6�׮�K�~��-��g�v�Ս]0fgVQ.��{U��yt.� � �w�v�h7u��R�9�?!�:M�=Q]k���ء��;��� �(�� LYP%k�|g=>J�ܳ�S�0�a��8>���p.��=�õ�#ůY����Z%6�F�Y#΂�Ne����<����u��S��L�nt����5�D}݂Șm��Ր��x�{a�r�ܿ�V�x�ᖅ/�v�J�]����h���bz{�Ҿ��E����
o/i��������H���k�;�}Иn�Z�oN�����8Y6��9u��=�W��c�ly�ӎ<ǀr���3~0:^{��Pm���g��=����Q^XF�.W�����~��ǈk�+�aG�8֒}hkMT��s�w_�MI��m�VaQ)z+x7�Oo��Pl��q�O��W��6�ї�)|V����a=�l�Pva
��L�-q�#��)�{R0\�@y�Yb�0x�u�E�/�i�#i�|�k�b��tJI%�RC�?w�^Xn8��|*������'�-�?�e�9<�fR$4�V����<������y �Q�%@�q�Y�'�k�d�W64[<����ɡM�eȺ|�r�E��V��W>%e���y�:yczcF4�����.j}������n�31}5�,�X�d#���
�!P���+o����ہt_:音=�]68E��ˌ()�������<Fw�^�8.o�5��:7ݙ������K���LuV�_@x�����{��M��aj��⮶��m�2_lG]�)
�(��	�ˆ�alR��#r8�:S��%)?:s Ko|�60�m�۟-��w$��b�#:K�M�MIzs���BӡBߵ���=p?�N��`����� ���8H��j������~$IX�n�\<[���}U)CX�'��e}4T�Ua$��@��I��mo�M?�W�Ś����Wjn6'������IԄ��FX���f2�vY��>z=-C�ֿ�hH�I���;���P�:� ���n��Y���ys���7cx���t�E?/H<	�P=_M$)bR�����HC_J#wZX���SPJ㨚�a�v�!\t�"C�ѩ`�t���3.S��+��!�}1ݻ�m������lA�g����O��*Y��Vj.��M�I���P��R�;�hv��a�f���qC@9[�3����?_�����)�O�B���2�-�b{��V:��P�g��a������� 	��"��7�F�ﵣ%���_��%-�</�s��X�әU����K �����8���A�J�Ջ%6j��T�R;�]���}�겂�<*��[��I��sk�U 2z��v�7G�q%H;��(	V��K:}zEtRoo��8y�;�Bi*�(I��g���w��/�]��~Bۖ�f�ҞD���G0=�&�[�.)u�"�.c� ^�����$�i��@j�M���)_KP0�gl\g���iEԶ���<��9q�w�R����'߶;��k�bt>T�y�|"Q��8�B��E]���9f�ze���4��V�)�#V�Ћa}b����(��.?|b����A�ɬ��ԑ�%r�
�(�lUGR/�E9��.ٚ��y��`LdfNE�`��>��RV�>�U�M�p��M�X<�j �Y�)���6���o�&�0#J��F�MS�eE��K����4.�g|"099y���%[I�RY1";u�'�}ݬOW��nʤ#��})6���,��V���>S�K.�k��Зn��􆧚q^��.sX�qFb��p��~L9R��3H����k|�m�<�N҇j�jSw�l��Y�:��-!�gn�����m��E��_hL�Q?Nv,�k�M�!���]��=JT�w�?~����~�Ѝ�dy��*_�����2��v��-t���Cw���V>��R�^�a(VD�4�Z��]H`@23�p=�v\I��
�._��JܸW���γ)�����i���b\cLL�P�m�����=9��X�
��E6v[me<)M@J�^��Q\�ѣ� ��~~���ZL��5�؂N�ϘN����-+<�b����l̢B�{�K�;)ʊ����|�ϗ�{{{ێr�!�h�u~t��1�.�9̖p�y�ISt�)y�Ҥ�ECc#2&��C�10��{�j�ڠ��_AW���rx�0~-PIF�L-ʊ���~ඨizL�J��O��߄y�e�~�|�ZDv��*�%�:n�Z=v�.�-Mb��!6=�ĥ��g�2��vٕ��v�����Z�U��T�E��^��gWl�{�J-�s�����"�Ss�,����ﰌ��mD��aiR{�����N�T���-$xת K��z�R�Я�_O�×	����XI��HF�y�=)Ob�
Q��UJy��<�*���G�N�K����Y����j7!�R����V��0�;v�x�R���T [�`���d.	���P�fj��]�c߭��?��,V���������,g�lҚ�(���˲
1�mé@)�'�:/tf��z��ݼ�������̃�qq+Þ���������(���j����{
R1s|m+��a� :�<f�Nuܮ����!�Df�"8���W���~'��a� 6�ˇ����~�+��B5�Y�u�nP��ľ���N���(����OjM�I�9G�@ny���&�`
)�j6N� bj���t�]|u�E�L~+M?�l�%'w�b�'@SRT̗� (�h����*���������;2 `����zj� * d�v�i11��:�u������'��6%%'�*�d��\X�Y)�S��V���~�\3���"���@0� ��mT�d)����;G��TTT�f{r�w(�>�<6���c�$�e-4�!��e�j�u����u�]�����Ri�-�����1---�E˿1��z!4�mj�>'��6� w�yH:|] B ��(����4��~'��;� %�u�
�	;�"�1򷳧�[�s
��iy{���B�ҕo�k-PY!O#��l �-H�2�ӵS�S@4q��an�KP%����2N� �̚��Ó!��7��Eށg]��3՜�Iq~υ�~ ��	X,�y�Ɨ���@����]v#�������_��� �}��J�j+z�}ez�ʂN�a/�$$�iX}�O�w����d�Ӣ�dM����r �Gc8��ٯ!��.�����_��	�Ċk<�Hŀ�7���5�%P��,�ɒ�~��nw�y,GQ�^f����ߎw1-mhԎ]�z��`@R*�Ĳ]�E�	8z�x�I�w��X�S���o�j�:�gg�n��o���
�6,�ˉ#�ހNr�~�E ����t�t�����U������\��"xSy���� ��q8������v7�����I�A
P�/��-���N�ϱƗ�rp�q ���#K� U�������m��{<d�o�h� ݪܴ�yW��~a�:d}> ��v��@p�5yZwY]��1�m44{�l��a���i�D
��ޞ����iu�҂���֌1�;��-d�
f��t��n�o�W��ٞ���)�)j��$��{ZZV����Q����Q�ee��s�v����ͽMH���אZ)0��s;�L�4��&�ᄄ7D��9�IK�����(Ah�7��HڏݎE8����}�^33775������	��V�����t�?���n��.J��`�1����� ��m(�ܞ������FUM(�{�!�x'KP�����k�#��~�T<��Ú6��F�d���~��	ĊW1*���Ħ���X(�.�HC)�E��c����\��8M��A5�w��FgO=��dTP��6m�2���/(n4]�����LI鴨	�U��&�]BA9��ʏ:^�A�O������/�Q�8b+�vnJ��K�2���������2�Sɡ��8�BP ��2�#0� /��h��j��>���SIzJe��՘fh����/���اW��z�"���N�+��?C�+�m��b�9 ED7�G�H\��(�6F��7�ܦ�����v�C�Pi��|�d s-��a�r�E�C�\��ֻO]�����/d���n<謥���*����K�$e����Z��%\���6AqǾq�G!t�!��yw�	�|�Wfd�S�<��9q+4�N���f�MFW�G�:�?�T�}k��u{�4�8'��� ����J�&
&�=ؕ`��9yy���S�n@A����G�Sz���8G�Yo�ԫf�h��@��h�kV=��_��UH�'��r�H��I�s<k�lKb�:��	��(V��CG��b� ������k5X��J9�?����JA� �*~@U��0.{�0{4�}�h2)Z+��t�ڻ�C��淎�yQ�2���p5p#��h�����ڞ�.�Az��
�#$��j�`ٮ�DC�+�޲�v9%�<�H��S���Cϡ��8-��Ժ�U2�nh���e��
+�P�9 �@�߃Hw ��{�@�����d�׾s gM��R @&� �A�nfvncc���!�)�]�����B����xf�Ũ)T#nGq��)�:zX�[Q��η��s���x^FFF� <�B�y�j�uc��^�����`�ߏ��u�W�X�S#E}��4G�>4feʧ]'=�����fv��q���2 �����r:�
�������@��2#�p9�W��C��@�wx�⏸ot�B9�ͣ��}�[�P����d�V?($1�Z��ʖR����p�ii��ܦ�2�g:��`�F,�ɪr�O�Rq��7�Z����9;(*� �5�-]ޑP��Pf��>"Pu�-4""BY [������8�TB���Y4��|h�֮���ܮ	��Šѭ�:z�ijiힽ���bfީ�mM���+�r��kK��T��A�y����J��zKo�R}�^^.��]�NS���O������F��*���f(�� ,��9f׿%<� �VXq��2.�M��^%F�-F�k��q� ܍K�t|���S���q=#ʉ5e����h�*����p�w�d[�-B�$	<���w�j��:�m_]cȟ�4uɱM1vhҘ:Ek������L5N��8�CqL뾄�ⓢ--�X%�`׻/ْ.���,�����S���`�ssj5���T3h����@_d��r1��'���/Z���Ũ�S��ܵ>��r������D3��]ŭd�����rp�n�S����"bg�h�U8ݮ�͒` �*/kl7 �_���7ٿ8N�����H|��:��Y��<p�E�h��Q�}���<�)O)����f���/��W�rpqz��芦|�f ��M�_�e#�s���0=p9�ec�4�<��H��}	C��nv�ck�@��;��8��- ����Ui: 3�|�hi5cLķuw�̓G�@xe��9 N3�H�.]���/���Y�?�H� ��p��Z�IEx�Z�0-?~��������a���i��1�?�D��WK�b�+7
[]{�f`N�����r2e��!�/��P�w�Ö'v8�5}[>tmt�V�i�ss(�x�N�|u���/�"5����#�u�N%��;���Ϝ����`iD;?�t�d������Rk{&U"����{���TP�k��[<����^������D����lJ����'Ų�Ϋ$�y
�U|�H�M���.V_�,B��.[H�s��X�l����g�6�����q�'��`aM���?U��ۊk߮<U7^ih�'�Ғ�0�p��_=R�kz���x�"��Qtn���ץ� r!̟M�[ګ�2�Cc����"z��������W�/ˌ"4o�ꗾ��]��&���k6겭�}�@��,�@��Sd�4��8�����m��zM�Ym2u����9����>��������Wer�Z�I�T��/�V�f��7i�C�-qdKf(m�j��0wf>���-�sಜQ)]w�.�Ħ����t{5�k_����Z��R��;�8�j{{Q�W}���a���ո����&{ٛ�`u>j��R��$����FX�����B�\9!O�?GW�V�g$�Ό%�oW�7�M����V&�_���P��A�窹�KWsf���K֤�p{�-�$
I��7����Pd��_�g^�J�\c���|ܒ��#�	'���+�B�0�}z\�*(D�m���nSg*�KǿMn�h��4t�����Z��yL>U����+�1�zx��uS�ZQ�!���Bq25�@!��v�>Fjj�� �5|L��mT���J�[O�' diҤxQN��\<�̙��E�G��q��������V�Ul���/y-�3���(Mk�Lq�M�G��yjx�s4�D�J���P^���@&�ңfF�މ~�s�����sJ�ǂ�mmtL��#�褠K�H���W�=����e�]�&$W_�����R&�ۑ���%�q�N(@z;&�`�3�[��n�3>��I���An�����VBԭ���S�#���j���}y�2���Ѭ}R�@;-_L��/���K�סg���{R&�?����DFW�p�����-r�E�5N7��'����\F�	���~cܒ妮�H:��k��s?�}�+1�<Y`��*�[��^�?0�X~i۲���)��>�]��������7�%h��r@��d����jbέΥ+G��[�o�_ q]���Cȁ�������!�QZ�pi�������Դe�Կ;u�+3�Wዑ}��ܥ�B�p����fmog��d��|���v���c!W�
��[��ǣ�"�Cy��ff�)������h����J�ϥ�#�[R)1)lpq8Gu)s-9v4 Y_��l�xj>p�Le�1���Ӽ(���EֆS�&��Xڵ�B(��kے<�e�cM�cw�X=<�5�S첤��Ի�bn�����O���l�)\���0ԨR�LگC���"�/) O�p_-���|�.aHnً]4�a�{�7x�D	�xb�܌���� �)��R��d�I궃R�B	��>PF��Z_^|3���������'*W�8e�h2�@����F�����te��/�{�}Ie�4eU�v��mll,3.��]fI֔�R�b\>ݭ��$x%ELJ��[-læ��+�HI�-���34�f����=S��Q5�QS��twN�sc���~tl�������7�N��4����N�u4���z������T�����^����;ȁM�`wc�k�m-�mx�&1�����Q����35����2���b���JA�� Cp[[*�T;|��4py;j_l�o}��b��B���e'�������)ug(y�l|o�[uOᩀ�[c,�rB�kn�/�O��i����%�G%j1�}������������L�%]�!9WB����5?_W͛���}ɺ���R2�;7����P�©�h��R��9�b����^ܤS��@�A��8�fi<,]����XNv�Y𝿐O)������P�	nA��LW��[�uF��ud��W����\p�"��� �G.'\�,&)3�ť�U��	O�隭�W3W|��!��q'�SiZj�0�d.��(Q@�J=X�+��lP���5�
\�u�#��ta�Tfwi(/��R����v�K8�b`�9�@�_��Y��z����E��������7�ٝ9Z=�m�bśT��#k�7��3V��XY}Y*�j,e�Rڏ�plC�����]����>���z���Pk�x��t::��b�ht�\_Q]	!���d��{Q^�����[O|^D��`����ތ��\<L�/��c�L�Zx���T5K��+#����Yg5�ð�F�&��=��.��%����וڛDb��]���9��6A!k[�KF�������aכc��[�q}��	=j��E"��aN˼+����y�D^��+J:��D"
��F6f�A�1�2��E�Ǻ%0`���FT�/��P&�]g�F-F
���fL+����}�����J���)��6B��ySݞ��,���*�0D�E�uԈ�r293���m)R���̠�3���>E}�H�N4ǘZY	w�����30C?����%�b��������i`���	;M~s�ŭ�g�Z�ϟ��4��Ͻ�_tp.ɿ���'���6vI�n��<�+��v�ߝ`��;�+�A�l�纇?�f�N	�K1+���;���q�^cZB�= ��k��Qʂ5*F�!km6>�t�\�Zy�6	���`��۾�����繐R��W&A��VT��2��w��c��b�2�m����ks#��wV��x�M��`�'Rja8e�@�W�����Ny�-xY����y8�,!�L��uj�8,'��uL��B>�^�Ⱥ�!�/�d��?����Ny�0,�5P���@��`P�������> }�=iǌ�uIS$RP�~Q�n�G��s$'�n<pxOE��R�$7�h�8��4Z5CV�Sjҍ����.���i��^�3�~�k�6k����Kͷ�y޸��@2WV�|��9�g���$
�s+��_%e��o͚�Te�
_����
�j_�Mzgm�>#"PwCn�=�|r���d���x�8�䳸K�A�=�oXVȊTn.R�(��~�lՙUd�/-��mYl:&Rlҙ�(=�*4H�#Q<�w��J�փVj�7�EQz��%$u=���]���Tn�U��Ў��������Z0���b��[[qLW��b���vB�<0�^��tUx��GX��������4T�@fm�%�)����ׯ7�z]����^}4Z`7�D�q"ı�;���@�q�E�2�p~\?cz3Y���w &��0vJ����EZ�Jy2?����6�}��K�F����Z]K����ʛ��638#�l��/ij7�c�כ�(��
'��V��q��G��t�m�̨���?����b��$Y��9>(�,k�����}>J�e01�/��w�V��3�֧Wߧ���-��;uɖd(�2�I!�N
{;Vq��%i::_#�⸲x�{���~�z]@
^�B��l���� VOB�nm�����l�ş�)�u�W>KG�
��)䭪����n-⤭>���
�B�~�
��#�B��E��A�������cXK����S��Myt�:I���*��|;�Ⱦ�~�P��5o�=3�_�<14���X�j�N�n�fӐ�8[ t�L���_r�3��b\
c�Vb-Z	�1'Q��J�x�d닕�־ZR)��C�u:H��/8 ��2x�Q�5w[�t3O;j���Lc۪�C�3�k��VW�+��C��X���ӂ�����G��F�͊n�O �[�q5��w㽉�%,D�س;�0�"D���S���ovt?�3��şj�e\��_�D�i�Z�#��e�����~��bR�k);�������{ G�!"ͥ��ovQ
h������Y6�	I�{�T��w"(�}ޑ�
I�b��a�[[`��@�����8�|�z�l���>A��XoԌd6'$��R��gx�bNp���[�q�Nh��<��A#��3�,��=��u�^t�yFY��40�S��Sq�렌��E&>�Ĥoԍjiűa"��'���Y�#�^^���uY����0������6�l�%or���y<�!�ln�n�,�gW+�m�n&Y~N�R�b*ێ��|�ہ+�<U��N;��)X!i!���_��Y� �$��&���.J~��n�+���]�ܿ1�cNx9+�D	܉�T���O�8������_��c��b�=����s�9��G1�����֣��JO�����3Z�P}'��Z�S}��cr��䁉�/l�o����t����Α+�mY�R����٧�����,��[�SG��+�R��[y�� l^��.uvypm]�x�A����{�?:���l"@~gI~ga����n�o�p=���*m˸��L*�������B�Y	\A<����8��"��^���\�0�_�8������I<�n��|'�I~k�L?�VQtron�1bK?GzX+��r��ÇP���^�!�ԝg��[��7���C��Ҷh%�ytE��te��qU��v]bRX�d��kv.���y�ܲ�s��cW�E?�</��!����ӊ�;�4G����u��nѼ��͆2��E�5y�N��ݪ��T��]���U5�����<9�CO��I�SYd8��^1��G;b<��zfk�fk��7���fY����F��g��r�zK��愓���+��'�.��,���,����Id����uu������D�(�B*���~FcF5[�h�-aΦHіԔx)���(NS��;�q�D �CS�aY�����;�esVO��L�`a��,�-ϝ;��2�a���a��i�ˆ�Mdӎ1���T��TL�O������9�9<��S�ɒ�降��q(��7������VZ�b��.�����y�= ��-�����bG��Q�6J��F�����L�=���R������X]���#1
5�z36܍���U�ny0�,��Ef� �����P8e6����,z���!A�+j�o>�e��C����B�̚�g��|�@m���^��������xL5ή��A2KN%�G�����d��EE����`�6�Ʈ��ў����z���E��%"�����:	̿�aeBE���E��X��S�b��:����EǱx?z9��P�O�E>�ϩBNƺy(mKN�l�#у����><�w
P�fU����,��[��77��ѯ�${u��)zM�F���Λ�e����U��G֞��=y��'qm�G��j�1|��ݠJ)ʃw��=�[AW���A��TU夂���[�.�eơ�}�zJ9�+mQN�Y�U�ם.e��O&G��ŭ�Q�4Yxܩ���L�V�K1)������I�����,��'8VF/2�!I�z�Y�����;L��`�L)b�D�w!�pH!'?u��'w�ɕ��-ɯ�yI���q�b����W�C�~��6�I���e5��z1��֕gq>���Ք�:�d$�7S��}s��2b��u�F�p=J���md{�LA �`7ZI�<(��� �H(z�E��j�����[dWQ�ѣ��$`�0NS)@��Z��`�ԕ�u{�6|.�ol�LI��JM"��-]�_�m�'����	���n[d `@8-�*����-���`ƶ6�pf��"`0�������?�7��є�sQ!y�+��KeOi�lr4��cX�3#���Kfs�j�tė��ڃ���z���&pO�r%�}�.���󐎽o"��<<P!qJx���[z�RS�^�U.f�'</f�oq�56Gu���\�R�nvN���_�7��a�q�������\��b�ݳ��L^9���ᩇ��~x���!�W�ttI\��?�z��6��/tO��TM�;���G�6�Y�ҳ�9
��D��O�����@��_	39�����%���%��7	V�?�_ �?��$����T�'�bމ@���%��7V��̂��(��������@��������+t}�IHHD��:�}�������:��0���:dc� ^����A[�g{C�+�n�T�����5�L8��r^m��*��.�DcV�OL/�K?'�z�l�?�3�yl�������5�����ݠ}����t����x��H�[+�*B�bT��ߑ�_t��N
	B\Sh��g)"�)����Z>Wd�4f���>�m�j����318zd'B�%��ܞ���W��-�vE�^�m����)���ĵ�L,�Z�30�W���U����[7����������P����е?E�Q�\q�_�ɑ#�j4�W 3��@����ϴ����9�Uֆc9e� ��;ۄO��c��v}�����Q���o���,kY�M>	?��`%;��y
P?��gg��x���(���7gnK7�t!�� l��J�=˔�VM׉�6�^�M�ߤcd�7���=�7����|GHdJf�p4)p���]�* �y'�V�'i������URQǎ+�U(�Wg���A[������9�}��y�v�c��g/��!����o>�m��㧍�$�k�kM�'n�m+l`&�E�=�e���o�1a�hi�
;��,��K�m�߷��+�ݤ-�P�_Q�\���W�AX�.������H46�x �{G�6�#����l��\��kS�~�[�� �m�q4�%��+��$����,ƙ�[�+�WW�=���g�-�r��A{�W�W��_ �24��ĹW:�����}�&赯�݊o�f��u�{����0��j�l���c�V�m�v�����ـ�7�e��B{{{�~����#(�l�o9x����ݰ����{FK����j_�҉�f�s���j�V!�J�wre��reӗt��f��3t���D|L���4����/�
��V���mJp GPh�� �y�����b���G�����cM�i�=� ,�`υ�F�hj"�B��?�V�ޮ�H��Č����Ə�)q�.��p�.�S?a~m_�S��\2���lZ".�/��=~�͗����9!�n��8œ��u��1ѯ��M,.�G���l�Udm�?��{�����oj���Ɔ�0aV��]aV�V��g�)�s#/1t��DG�yQ���`���F���Ƃ�y�� �֯�+�W�j��r>���@D�R�2���c�j�{�x��V��/�4T�bu��6l�JT�8��Bx�D<�F����1237?�^	���;�>��z`>�j�	�δY�4����5�m!Ci1��F�yЇ��V{�����6����p"�c/e}I����n�G��bݏ�V���z[ܯ�'�9l��7G��:r@�6�|���̇���\�&.�k�Q!_���rsm���؞VFdwyQ�lA'�qK��*�cam4�p2a����G��6���'M�ϙ���?:D�*n��g���ŗ��Ro��X_^
����xnO��Z�-"S��#��׬�r�zT���X�d�$�x�}�����KoS�,dm�����D�x��t�┬����D���1�7YK��GP�V ;�����vu�8v���$W�4b�� ���D�|�ul ��JN��4�͝�%��Vs��p�n���mZ��7I��ˀ��.�&̺��W���m��H�X���J\c9�0vH�MM���r����\���1ă��&�ܢ���ty,T}����ܥy�CWt�M�l{{�z0�zp¤!��u��CĤ�X>��b�`n<=�AB�ki�5}6�=u~�V�7�"�t�m�p����[���=e����&og�V��/�p�ז�3b��(��X�E�e�6�Jǔh��m|.hXr:U�HPml^�"n�B��I����X�`��N&6���,��_�޴�A����a�4r�.4�/���>��%�����L�|��5#ٺԶ��oG�d�EM��U{��������=&�?�y����/C1�ĿԶl�X��FY-�?��ŞjD���J.�=��g!��i4p�q�%堪�\�k�]b�#C�_��t鷓�>���*q'{����%#��^�j�p�ޞH	<z�/�8.����l9�'_�Q5��Q2l~ظ�ͰMS�Q����u�������F��C�6�������܇U� a=��O��͖Pf=fդY�>}?+C|�p��X��Y|�x����7bw�ׯw��K�.1���'�vUt�I��bTcUA���(�Bv�,��3Y]b���>Ԍ�x��Q���v]�a_}�q�p����U{��q|�ك��ǸMu.we�/�浜72̵��2k�'�&,y���v4��Z7De*�����b㔸�Ƹ%;lBq�P��ٵ�N#�O1K]/��vA<�)`<���G�L�8g
`oQ�:�?�p~�Qcx������Rx��M�cڪ��~��u2�y�O�|؝;� ���wF�u��<]�������s�7V2���a`e��U LL,6۸#��S�SSSV}��+�Y@���{p����ߛ
"u
��R����_��qȼ�^y3Qh��
�HNE'�w�þa��x7�R�B+%�bu1)��O8������b6��۞[�0��z)u�bOO����gb��HM�o�;����U4^%���8l0ף�g?��x�:��1K-�|{r�e)	�+op=n,	�yV�(�*�֍��Y�r���sz��7��Y��A�57����>�o�D�aм������֙Z^�%l�Ͻ!����t@J/�5s�R��݉]Qy�f!�j��)����G��楀�P�v��AT�c����]F�����*K�V[ .*�դ���'�k��b�~Rғ�Vpb�ˇ��kMV��4���ҿ`��WM��W���Ɵg�k*�]�=��43S�t��!�<f"�K�ؿB�V�7�X����o��6��Z������=D|�:d�%�_ߥ�Bm<c_p����ۚw܁@��3�@��~�ǟ�5��.I���$ޤ�D��R{����r	zx��J�z~���y�nLtKWjZ�Iu�2�G엣��,�E�1@:W�2�e�B�� �TZ���p}�t���I��;gk.��Z'�w��\tqG6�n>4������Y قș������#�1�~|:O�i: �U�c�A�!\���M���.sO��f�}q�&*v�� ���/�5Im��Ffl}�ٚ�_To��ӼR���'������\J�Y76��~�<��m}XʥC{5  ����mԤ�+����]�]�Ƶh�H2W���Pf&�I�g'a���"������-n���M�R��`� {����8�����Y@�Q�O�w.��x�$����7��ЉcK�S���	"�n�_g9C�F,���Aπ��G���0�'K�V���sA]���Pg!���4NG�>5q�L]��H��}�w+��>.Ԭ����xB���^�BW�U� J�U���h �ۆ~GI���8Z��P8�m�ץ�)E��G�ڞ5M�א���ęC�K/t_����Ԡ[��Nj�*�w[�aI^~�@��e�h�=�NMݲ�=�b�JϽ L�Q�3]�$d ����E�v���"��#���R׫�7�Dj� E"�������u)��Bw���Љ9ð1!�;�?��4to�a�����X��	H��]�փ>�µ�50�"�}��E.]9D�&��1Us��n�jІ�D�Xm��7��بǷ��[��7)M���D�Yl�.J?�a�q�ٯ�]H�����J�SV|������	sUe�(w�&N�^��j��1�g����ɪ|�wƛW�7g���i��1>�]��C���O:ޣ�R��*��P;�=&m�rn���0���w�p��#Zi`��.�ׂ�W��S�*�6���u��y2����ET����Ε�5DU�k�.�>��NdAI���wΉ���Q|�`�z������V>��1������M�Xlg�.��F���5#�X�N�H���ȓ��3�d�#�4�16�t�����n��U�����!��S˯Z��P���n
��(�+�߉��f�:�f5�\I���>d�*�Ib���Nׄ�����SY�TA~����0����̢f�l��NH�ӧ���v��H�q���TZ�w(�?�E�o�O,��tXo�ay"��aL"�?���9���!LO.Ht��Y&�|����M}W��p��T>�m{-e��ǥW�Dͯ����:镅C�����x0?���jML&J.7���cU����%���3�i���$_{�M3�M.���ۋ�|q��� MQS���M��x�k1������"ቡ�5~�G@���?8�JCB���6����%�.��A<��$Kh�^���y�ܼ�/��{���~���Cr6���v�w#�q����^瓜:K���]Ľ��	�����qM�sE<�u�?�j�Y�h��E�̷�n��%5�p�YnE^[n��3�����ƺC���O�!��-N������譡��a�f�"w��L�ݥ��,f���a�.����i"�-����l�������EK�ʃH��;u����N>}�F�B� ���jHX~���=y>�n>V���{ay���l,bMϢ�_���7dt��x��26ͧ^0pS 6��5�w:�g�c�(��kn��6)�x���3FFN�F濧����~�����"+�� ��]������e$�k���?��&�1����5Ɵ�:�7�*2����p_��QS���/h����Q��>U�b)�6ݶi�:�4��h��S�Rҕ`����бe���R�	�c6ӏ�z�o��gy���%��R^�+�А���♅�]��Į�.:3*l�H�ם���4��·�|>T���T�+QL]F���q<_}8EV;�]�b+0>ouqq/d+$6~�, �)�`I�@^��޳|�*l��v��d�`_��@\�sl�����WjeR�.���{I�(�%��V��N�BvB�̜c���C�v6���W�y8�C�?���#4����QO���2s)����k>c��Nԣ�%R��;���s���|o�֣��Ӆ�|5���gG!�������^%��*l�S^dɟIg�u���O�G՛#tN�.z��M��8���5��i����ό���y�ȥ�U��,>̀P�7�Ɵ$�[��n�
�0�*OM�5��r��ta���7�rZ��@W� ��Kw�z�DU�g�&�'���v5�Kd�E&= �! �dk��+]a��⏲�W�녇�t4�~���+�3��j�Vr��9�LC���Q�	)t��L����(K��T�w��/�Ԇl:͍sfҹe��E�WK{�BB7����*-���e&��'MԱO�ؚ��x�B��鉲��"�K�k������MK.=��p1���y�=����PH|hr�b,^��Ϲ�w��l�b�f6�<z�Oʽ��қB��$�Df�7�p/�|��s�;U�1���7h^��V4��?K㈿�������N�D�{��)�����_�5���o-_#O��SÕD�c�~hg�䢸�O���J��>��`���|z�� ,G6�iɵ����pa!,���P�LOJU6�������j��!�����&�,Dw�`�N�YE��W���w	�d���'j7oa���0A.�coKl�����b��[^qtc�k�@��LM��'�o���P��	�;���Gl:`����(I�e@)(O�]iB �q�W�>���K%�*�6t�~]��k�ub� ��;�����N|:�침��{�oU����'<q�$�T>�����ys��N�R
!}4��-t���Ѵ�
h�?�e6g��Z���ӫ�g1[���.B�B1��3|UFf#Dڋ�by<�K��B�?�W���3����d�M�����3a�	~�o�!w xh;�na��Ĵ��A�Q���)%�#W�`&Uǿn&�D��������MvN�R�U���G���Ն{��9!!K3�Wϟ��8�~̲{B^`}���j�k�d��>��R��?���y��Y%>Xq���pGy�j��I'S��Cg�*��D�k��=ZP7���L��\�^m��p��UH�%>D����$�������<~���#t,��U������M�	�$�B%�7L�p�5�����J_=pz�� 0����/��iĊ�W�v^R���,�nt+�A�Y����-�%��g���-�x��vt4z����[�~�����Z٘���2 E�*ݴ���o����L3�M�*J�և�ɠ��R�8�9Z���� ����Ak�����P_{Io�^	>�v�p'X�����������]n���m�L]�̤Ȭ�!�(SfJ����1��2���)���2Oq8���1��]�v?���=���Z��z=_�����k�j:\Tأ^/v����uE����R� }G^+il��>ɀ-,��su�nl���R�ŏO;+�[��[ ��D4�������s�8z{-8賡a�/�>���~
x��$?�7
NF�rg�m�B6�=�iz���Ʃ�����眵�KtZ
���:E����O5=�dm'(p]*�H���B����ss�V��E�9��>H�A�H_x���I�s�}�m�Sfqc6��/o����C�p���J�u�����=���/8[�_��-���P`>�iKp���ε"�y���`6!���e|J{z�ʂ��p�ιy~a /!]���7�[�c"e�/6���(���?����Ǩļ$��-��+2DL�u3P�
ޡ�/Q���z@Cu�V�iH��8�P�{X$Tۮ��?uj��^ps��[WDO^*��nN����%��C�gdt�g"��/��xC��E��%��B��S����ŵ�z$C�b����0eu�9��\t<����5�=g2���+�5�/��3��e�9['a5�G9���7�뀩��.ǧ �O��]2�هac���8h<��8��腂-{���.�=6%r�oo*��"�2;�C���E�J���Yl��6
K&�;`�=���f�4�9kE�=��}��>�rO���}�<���	�R�{AD��e%�H\fy"��ۄw�f�i
�E�梔�tv=���~����}�zd�^�i��}<d�5��kg��Q��j�=�{�P���0�6�1��lW� ����BH�3�����f�Z�>���s�%��\	�Ǖ�LOd��ٞ���p�{J|ieI���5p��Ԋג�UU"�:F#�n��쑛��[?��'� X�**�p�O잷m�z�lA�k5�D/
T�/J$�+(�P�J��Zy��'_v�fХg
�cQp�^챙"�^{]��4Z{IDi�t�{�^����uD�v;����K he��B��k�(3��O���}�Xk�[�wZ0�(���[N���t��9����4?WT�x�7��E3��)�tW�_^�$-~/�����U@;B8�����ʵيhx܊����,�kU�������mω��, g~��lf��"Ҹw ���,l�QT
�$z�~��r�.$P^ ����߼��U�C��\��ֿe�0ف��?��d:���&�m�`2hǯ`*�⬿oL�!ꣲ�u����R�ZC�ݲU�v��Ր���@�\b8c�
��F�}�� �2�q"� `gO���$�y�#��y�=����q����:�8g�`�t�.t��B
Ȋ��S��4}�F1���6����HK�ٽ(W��W��c�)����n\�iȗq۬��ת���.�x��g(7���?./=o���b��)�y���R�bL�	�ѡn�۟���kfC�~�'��S#��p+Ng��Õ}���z�I9��?��^��U�2�m���1P���=Z�a�l�	�:��>�Qt_�G����P_��[�Z:��ON���qe��G�p�^ n���\�9R�]Gmi�V�ȯ.+�ߡ�������V��
@ș�w~񫋂�5�����{�G3���c���{���V��/WdB���wVQ����"�h ǭ[Ğ�zY���(�u8S">E(n[fɷ���Gr���B���aZ)H�N+6r�R:"�e�F� �W	u�Q����S�6�V_H�?j�|��{V-(N����(��:�|�\w0��Z}]ۺ�{����#�a��ur���z�	��W��4�7�)�4��B� \j�Wj��7^������J�θ�<�7���x���p���V�>���.?��u�
G�2놧��!��;��C���+�ƕt�3ٝ]���
ؒMk�3�_�M����)pq���Z��E�U�{	ɑ����Ķ)����dm5��h�-Lz_L��b�(���/N+��+f؂V<J����t��u��@/9j�DWg�����%&��D4�w���V����t�1�l����A�ج]���S� C��)���(�bUT0:�?�
@[��+�8���e��3uG��u�6t=�_���N@��^?V2�PI/!�v��0hX���솘��<��>gJ$��h�����eFھ�%!�G�&��R��/嬝�C��O��4/|G#m����i�&�f�D��^o�=�A��ske�c9�Iolǣx���{jq�=���9o��\�����'�,l|%��� �[�@��$y�������L��E[c�L	�;W{Z1䱃H���3DM��i4��1(�G�bhf��
��x��x�� \'s� ���G��Y�D�H5����G���Wq��#���"�#їP_�d����7� �d��X��:�~t���p���E\�ФsxFF}th�$8���7��7�e��:�Yw�� ������f`�&	�˷;`o2OF��X��� -��8�}�$)���O*�H@��HM�Ϙ�J��Ģ�w ��:[f��E�����^�HU�z��0����9B1�S�T�#LLv�{�U�lRT�#$�(7}�u+���C��N�Խ��B�b0]��JC~�M�C޺��t���Ǫ�[�#㵊��ď�3�(����S�ſ��eS`F�hҹ"����e�Ѽp������(
���	W�*1��v�`�gR�X�������?��� z���gT���L?֘��T��m��B۞��v���9G��]읠�5dzFd���`�������͚@[QB�g������A���M�a�#��"!�P@���ܜI��dQ\x�F��.�f�dC�J��P����]��
�m�����������;�.���iq�yQf���15@5[c�rqT�hх˙��J��c���t]����M��w��>���\�-� ����~��n���`���E\�*S *^�6��-���:u�L'X$)�ג����}�K�q�;/���/�
��"<�yzgBbz{�=S�E��itz�[���V1�r�U�2�7�1��:�΋`�P��b9;��[��Q�<�Z^��9M�vu\]�:���W2�]5U�i����t�������	�؃P���)<��`ke�m yF�K�s �_�멿�\�c�t�n����)��vE��??��`�ǵ���ygi<^M����;�~7��)�%���9&��MpI��,ՃH0���gw�:����'��ǟ��S5,���sTM'�61�-D���q��Rcop��kQ�
FwzT0=!�v:'y{$����Դ��w�=��V��ơE�����^����_��U�c�*e�m	-ά��D����m�TI�cO�����n�	ܿ|�ǂ�b��q��s���l�ڴ�Z��q_��EH�.O&����v���w�4��7Z
f��D�l�#/���}N�ٮ�U�:����=9���-H� ��V&��_L�l74�����d;� ן�+\�5�9�]�¢��\�b��F�\�-U�1w�	��aDlʚ[��Ƿ|d*��i�����V�8��\'���y39~�@#�'fz�a��@� �aH��J��M���7��M2{���-\��70�����=������,�3I��nR7�I,�,zn|
�Pe�����/��:��ͧ{�VzI[Qwn�jG�Ʌ ����J]�"]��T���I��7�+<��(1D��\�D+�NG4�L�%^�o0U:�����P�������E���3�otB���@�9� �B(��жD?U��õ��`�gD��o#�d����0v\21����s�d3�����X+�QI;k8Bޜ&����ǳ����e��y�����Ƙ���vXl����E9���6�����va��7�=��2�Bv��Tߺ���/k��\(�����%�6)�u&���{{cv޿�P��x�o�_�(I��r��??Pz�[Nse��a���^��7��3|N�<� �g���!Iey�j��w�B�'Bb����ph��+�Nx@2�����,T����f`�����â�\��|8��JKi��n5qä���i���UT�CEa��4�]"lP��K��V��&S���r�����AY���7��I���	�1��)�|
K�����3�an�>��2��h�3���#�'!^��U���ij(��E��;�Laz�"ӳ��BQ�]���A�)5�L�s��T�Ls1	����m�%˘�N#����g����4~���(+8_t�V�\:uL�|2>�=�3��	ix��K���qm̔آK��;8)r��3�ͽ�M�~�\�'xF�̤E��A�+7�L��kU��sʠ�V�ߎ���{ul_,�]q 7�\�E�hZ�T^f߮���ʩ&��E�^�,�ߴ���S�f�ה�������>$�n���qgS�l�-��g����N|�}Șk߶�V�DsE�����*Ԫ���?2/�;��K��U��\jy��'U3��/o�o������:�&��R�\�RK���Mö�k�8�v����H�� ?T(rf����wiwU���[�TF�И&�9U����	*�����d�Qg�DXP���h�����DC͚���:te����3�ߓ���:v���󫮮�l�ט���:ԕ��u���8-�qӦ��@�4].��f|NĦ�*s8��Iz����:F��xDԔ�6���hb�$��5�9�P��b<e.�@��E�[uf4�*0
���s���i�(d|�w)�M�dwM2���W@)���?�#�e�ܭ��[�)6j���ޑ��a�rc��O�[uf������K�D޲ �e�}�ũwʫY�����!w.��teb�_mX�� Mb���W4�5�9"��֝gl]iۑ� ���A�)�^>G��Z��T6`� �zz���k��xv���Y�(�I<��d�fd�P6P�Qk�2/�y7%����:�:]��Q���ȹ��R_Q>�z�Ӱ�N�~�wJ��s�ߍwDT�6h[\���I��ҹɎ�r���m�ŖE���v���;�T)�X]S�]���vc����#6Jr��dȼ`u���G�j�gq�	�s�|�C���.ՓB��NS�EYt�IQ��!���K����q�(��W�s���I����7�j�7����������t���	�^���7��Ê��}�pG���)�X,w�$�����r�^Lt�pd��\�����ƙ��9$����̩�+�U����j�UD�x�0d��XU��g8Ը�0�����[ID�PL;�_G�#E��sS�bь�A����X����Sv� ]�����v~����wV1ErHk^���n����đyCMowJ7ݠdr�I���Y��§��Fwg�W$�jU�=��dJ��{C�4���}NQ�'�����i��ɚ�}�7����A�3K3p���e�L��c�_��z�0��UDG�ot�R�+q�f��$�~�T�����^0֒��g�A����rs�m��߱��w�����3{�
,n����P�"��L�l����>��t
qW���w�,Q��K"���Esi�h0�	EKE��p���韓��z
T��7��g�ly&Ip0v�_��Z�Q�jqn�7/± �9;����܆�O�[��K��&RHA%�wy�1���l�}�O0k_��'΋-���uE(��T����H3h�|�1#���ct�|˹N=&xփ\R4(�=��1�1@�())�P�gn���մY��0²��cPl�Fz�Q�v��}�fp���3�jȷ�+���7��l��f:N>ʭ�-#�HK٨[����?��a �WO�U�^���-~��w4	,[��&�>� .�P
㩅���L�����嶫T�T0��*K e}V[���"a�5;KjP��d FW���㒊����ʊ�Y�}� {�㻼$��(n�lw���%��C��c�ؠ\��p�h[^I욹HA�����R@�G���3��Ӏ�$�����okdP_x������ۊ�	�uF����ϩH��X�(���3.��sUvQvxq5K ?1Q�+�{I*����Gs���ec1��74���.�������^�MB��A��1�G���RI���ސ�َ݂�J$a�ݸ}C��~iT�͙��u_�Aش�hʆ��>XpndxRu2}��0�Z:��y�����L���Bx����z��*������#Ώ�F� fB��N����_����R�S[��J�DP�+�C�|c�!}wBz�']�zPV~_���K�:�AeX����*��}���?�+OIQ��=p*��
���Ƃ�f�B;P�k�����ϝ�����Ef�~e!��e���7
�������:���I���=*?5��ͻ��t'�#4���B
�go�l�>/*	G;���,y*�����ցf�7�[�� ��j=J�%V�b�=��ѧ�J�v3��1�7܀37H�Y���ɱ|���**8%%e���|9�[3PBd�spi�N������p�|@^cb���4&�36����Ow��磑V�&��4_T�L-���w��|u��&��~�h��^���UZz@�~'\,Ze�7/�^: �"!w���ja��ĲE��'^�����Ra�h��d�qʫ�1=�S��B*;9w&>����-�7�x������=xAv�l�3�_�א��:ǻ��X[��P�%LYǃ������r��Ie�������=��VlA��2���K����Q�M7����0�DWg��<��Qc��S�!�Y�߲��I�Y2���h+g�6�����E"���}�|Co]���"\l���l�5�����*�8A��gM�1����2G���_M�lp/�_�F��`�;�uU���~3�V%?��� ��dJ��6���c�N��n�ڜǣP�>��_��CD�n��-e^�tʹɠ�h���dĝ��גܖ>�#W��6����M�����FQ���_�ꮕ�M
�?|���� ����T�u��=s���|`�چ��V��v�������3�p2��W���V�$�Uy�E{�����l:�<��*Ɛ���(�A.~��WB��A�5j}ghY�~�1.���+�T_L��Z�l�O��خ�<��|�*BW݉�ο6e�8+-	R9pXy=�0��:������b�.[�OJ�脤zc��6����G���qB]�UNf�o��M���Ԑ�;6M������y!����$Ѝ�`�)%��5�a�?�:t���1�ѣ�I�q�#3�?�H�j�Ϫ����j�9���������ysq�5����aD\$��#��ɕh�V�.t�'�Y~�;R���S����c��T�r�P��{]s��������٧>"�?��|��v�ˡU+���n�Cԕ''���8ɁS�3A '�����d�c�P�A�s*���sm4U�V��K#��N������%w��:)L0F�oа4���F�Z��
P���L�U�M��s��ѓ#�O(�g26�6]&N0��I��5���?�!��6'?�nQ-�:,D���+��L_�X��VS��_���C�5E �؅B
��6�a�	�M7�McY7ak�Y�P���X�mˉ��K���%2vë��Нxi�0ߠ�|*_��(W�b�nm֦T�)�7�_Z��W"���x�D߁�,{=�H��?W|V�e��.'�=��y������YtuM\���/��r��Z�E�!�у��>�h�[�5��j3o�:ڋR�O"�l�uoZ���7��g&�rq¸!��|������Y�m����z��������omN7{Sk�r/�*T�r~�*+�J��?�~CW��������P�ʲo�Jw6�ɡԭGrzU�OH���/�M�h8����wL^�������V�^W��=�i�Q�g�q�7����h�՘EI���_��FN�L�^v}�J� ��%t ��a�aY�%-򦶬~��d4C�����x��5o��2Mϛ��Gf|V�M��������+�Z}|�}�����h���>��@��^�C���j���H/a�����<�#��S����m"S�)L�T��3�2O���A��;����rUUmЇ�*�F�/&�P��)TU��<n+:,���>�����Hj�1l��*>p�ĄD��ۚl=�q��2��K�-�y�E0���R�i�Hg ��>՞b�Y�ﶫ���iv��՝��\ѿ΄�Za��,#l >tt�g�̓�zXm�^����f�O����`O��z��A�R_o*�")Q��K��_VD`7�wO�����⎴��j����r�7|�Te��Ff�$�{�7E�X��s��I��ZuKҿ���Ę�.vb��T����:s���#W5[��ݔe�g�81�s������K�K�_�\�%$/jH�O��nΙf.��v�U+�N�����k_�,�]������U�k��/�c|VS|V}}��.�{v�rn�蚬zJ�f��5��԰��";�_	Z�>�H���n�b�<�;|*NӲ��1���@��L�RA�e�a���EjY6V	V�/:�G��*�"g�N���[�W����od��7�:���MI^`q��ԗo@��։M�5
km����2��0P̺
@�IZ0̶���>��l5A�U6����f�<g�8��t����M3s��ZԢ��6%ډ���ʜ���ֶf�����h-ee��/1���_K�vF�8�g����qڝY�p'�zWI5@� zR��eM�K>�T��P��t\��n�sz����%ܿ6����c���i���fO��q�������Ykn<I��@]��m���O�5u��A��Nrb�9��o�e�\t�Zm�x��u��Q!P��][bӃ��ٽ�\��2C��K��J�2;�./�	�f��+�,/[e�,[u���5k?�
��s�}6v$�|*�q��8��^jz�:��=��2���s���k���~�e_���yp�ҷ:��|�tb>�q'@?�NPp��-������T��h�	�g��K���y^P�D2F�}@p-�jOK��Fv������e��g�-]\U`��F��D8�<�1���z��v���u�̢hw^��M�B���:�i��y�-~/,B� ����L��Xޣ�~oc&:����q�s?ێ�q�h�8[ad�"�Cp
D#��x���d�H9�ʮ{�>W2�5���i���^��|
�/�
ְ8=��Kt�v�:rd߆O0|������W�:��#�AC� �tqG׿Q��g-"'[�����긵o�)����:y��S������ ��ܯ��������兼2��m�u�&B��D�$փ2F����!N&�qA����#�K�G����?V�j:���
�:��I�w�����Ȭ�b]0��>��M��??�̥����1��������R���c0ు���m�?����M8�8�ghlE�_�Ə�� AO��z��h�A���O���S�l�H�\��r���4�Cj�B�8�N�с�d\i��4��駔��&�RPo/e��t�XJH��Z,.��8�ԸË���SD7$v�L���X~&�8[N���s̛�#��s��p"�����8���<�FDD��Aj����g˼�saJ[_>�\8�Dj�Ճ�?~������������J$
���NV��w�?���*�(�äƛ7��;(p�?�'����]��W��]�4����U�p�Pp���^�^����ܿt����m]].�C��H�Qؚ��S�;���FH��.!�cpP�Р|)���t�
�gg�$]��K�Ŏ@�H�s@qʡ8�`	YW����5D���۝��ѕ��Α����B��N��O%��N.�445Uon�Ʋ�Щ�$4�������ǅv_��+.C�T�zA)6<��uu�5�ޢ��fU�]$��􋋋ٰ?SCH�� �+��P�/��W�9`��LS~!]���	P"p����k��-#=D�nz��ťW��5��� \܄�.�@6I�1��Z}�����Hc�2{2�WZW3��& � 1P	1J|�j�C�u[�;��@����]3�}��@��M`��o��ӝ�3M�D�C0�Ll��B�|����a��e3`��P�+�d�I��F�9����Sky�h�_�VG�J�b@�6���P|�0�Q9|�:a��]xZ�@H���}�7H���cmm�,BY=1�}o�9��ty�H$�;w���{+dI�Gi��m]������5��+���p^H��e��2b��쬬?DIm��-�t�=,j�f�J`6Ε�iݓ��b���\m����)+�����G�¿a�x��/��vBӄ�B��TPXHOj�V��=��ÇH)6���M����+ߺ�{��Sg�X*2��c:���jj��K�yS��Ǐ��_�jY���j1l�B4��n��ul�^�����4:������G
����}а��|�m�+?�]�?0���XtJ���3R���+��Gܿ)�hhj�K��(��3�3m�=@0i�jbb�+�A�O=Gy`�
�!��Qb\|�bG������O�<����
I�3}��
�"w�<�G�m�:l��>^��T��펙�|���&W��ɾXۏA[2��h4��RM�3^��\b�M�W��8�}����	��[�����<�Y/)$o0	��p�S�2�pLj(@F��$�l��Ҧ:v,���6��klj
��ӛoc����q�%C����BA�*���~On]x��YZ�~�f��i{���^�vs� ���h�&T�0�����w�=|��C�Q�iM�W��?2}�O2W�X^�G���������R?@�W�Y~5���Zd�PAMԑ���9�}?�h-�}cEk`������BC\{�Y���֩n]�A� ujr��Y�,oƴy�aIMZ�k
�Tq,{�P�	�+~+нl���l�(�����l�9��I��|$�w�@r9��m�_'�ꨧ3YW��<J���+����=]�}}��F���~�����a��	�\8z&&�ngN�N�)P3힚-���*�����ع����8�-�F-�빜Ej��6w�nі%�.
q^ӽ��������:����T �8f	�
[n�+���(���d<��m���K�����-�{X3f�82����T�[W��\�|��5�t��3�6���D5�_Yzz�������h�*�-5�8Ja��t%))I��Iz�W��o�ځ��{����S`d�>N�(U+M.��~|��U��Dr75y�P��!w�=G3�>6��Dl����}�cg$ �o;Ȭ�o}9[U�ƍ�-�#-��$�Mhp��:4�e{�	:7��'�(?��܄��%�E͊ڏ?��2�p�բ�<�9ML����F��^6��c"}|���RS^ZX�j��~A�b���J#F���l�qUS�O�mll4p~����� ua͕��s7��m���%����q�HY���3�ֿt瘛8����+X�>U��E״����g�j�A[��]䞣�[����y��`��V��H�C�i��A��#,F���z��W�,J�F�����Ề��:k��7n�8WfY�]�6}e{444t�������ޮ�q�aS�� �N/��.����ȷ�n��6��{l���3R�x�,h��u�P�Y����4��M�g��w���˿+��q��G"�^I����٘��c�^�)��f���A���P�R�hS�8��Ӈ�
�|1�ف�����1i�ò	6���=�Q��{�p�&���T���� +���F���l�L[��q��=w�v����ʰ֘�^^>�j8�=sʚ楯�oW�����~��`7���P���p.j�IF�(�<�z:�f��?TU�2^��K'+��<���e��Aq�����ZXI����{�(�~��_M���o��q�t�W"R�д�G��r���P�.)}� O���j	8��gce�WP0�X]Sc��\D�uez�&DI���fH�F��ٗQQ�e��|׆�Qt��?�c��8P���C�jum�H_6;7׾�H�ҥ���rM��R��!8���W��H��(�����ӞNߎU��)��*����O�	dڨϧ98n�G�Ke�`��1����� |X�F�yHH@�Vm$y����9pBd�o�)(!���s�y�x4��zxH�ٞ�C�)����"�	l헮W�����8͕X�i��c�U�%���(��h�9=��]������	�y*�6S�|d&�����A��A.���WD���?)�}�?��\'*����=�:�-wnR��ǟ�J����$>�= �v`���A@�+�)b��X䈷�wɫ��
7//�G�<||��zy����if���x��M�%,I3�b%����ͬE>Y%���Z��/(C��pۚ2
J�q�BWl�n��&�:�>a�Ɍe�i��9�}���� �r@���
����gzŁ��LR�VV�|��:LWA�*�v/�j0�+���Nc����8�o���r�S����qP�ִ��e�"��և~}�p�ɩ0�$�)�� V%�*)�
�+b�DV�HRt��	�g
��&�؁|$� .�E<��
pi�(�D3O7���..&�N6�X��<m�z^��׍vUi&�U��Sˬ���AQ���r���l�`��Fڗ@�O�
��,g���l2����
��9�*�j�IM`W�+�w#+���{��L43U��w7*�%��V�dYq���� 0���Y���p�豞�)�i11q#H��3���[W�2ɓxPR��s����S�{j�n��j�Ν����1W���	�q�	b�п{E��{�;�i�$���t3��[��Fku�Ť
N��H���٨`�uܸko���>�9E�)���A&�I,-�`
�z���r�>(��2�Eث
����rF�XܗZcx2E�cʛ_Y�� �6��5U�QZ΢�
����Z�,�:��p���i�p�:��$�W�����H�u�LYm/��1�4��+fH��6QP ���2�\[��hXP:ʛr��[f�&i�-�����*��Gq��.i�B���(Y��O-6K�x��{v�F���j
��]��g�Μy����4�7xFd���?((<о��z�ʝ�Ov�8=2����Y<�s��q��@�4s2��6~�+0;�Ñ��}JO�"��:��@a϶�5���er�.+�qG����\����é
\�������"��G4R�t��ߺJU\��Q����";'�7��]!		Ɛ��#"�7D�O �O�c6n3T��b�kmW�þ����ʩ�X��n��nsq��A����{Dr�YUa, (H!Ow�>`u�^����w�d(wA� G�{��;�Z[[i�͒ѮI4�^=+��Z+-�{`�.�;o�B��+�azh_�h6��jO�CQ77�z���_(4�ū��;7g����� �T�t8e�<H�]@��q�Cũ�����fgg6�/J�,jkk�w��1��ǯQJӃ�4�D>�7��eh���%b��o�h�RK���t����"[��E�VZf�R��CUu��c:S���ty�]�e6L�U��R�jM��`ߊ��ȈM��/4�Ȗy��V�W���%|	�e�)+�	F�L���E��E1M����Sy��l9ŵ�+ֿ8��8�b�%`���O��4E����^��������0���� ��:���͕(�U�^�ZO�.eRv���p���T8��#eU�r�aאpK�\a�3x�S���,�)�;4���$�:�ye�����i�#���߹����HQv�u[���~�����=�<|\��g�c�E�P��,���R$�4g��V.l���1����G��F��{�O� >J'}��W A8<�L�z6�Zr#�Y]�_��s-�4׿���������֜�?��J%G���{P��E[ME (�Z�G�Ib��c�^ށ}�,
К���ͷ�B��\�Ə�r� �fcc���oS���ވB����eC��� ���*��4Ѫ��+ߵ�Le#;lq�6P��48�HhӁ��i� �cy������Cp���h:���7�(W��?J �1�;V��Yafd��(jQ:�e��x[N@�,�k?����s5ˍ�pC��i!�w  �Y��tog�(�I���>lS���&����l��
����V����2K{����C
�_�x�m�4777����<q��ի�S}���Ĩ=�O��:�)Ж^�>�_&��)6�RSTV��-9O��y�}���|)��h'��4;�w�@�v�[3&�&&q��8��Lh�u1��-��-����n5)4��𭷀+=�/�*
N�j���:�Jԕ�L�#����5�B�_���n���N%����Eח��th�o���YҦ5AmM5�d�\�{B�E�kK��90�9��B'�&���#u���ᗫ��Wb�j���B�Cň��R�C��SU�w�.�'�d��M��TWWGv&3���f1M��$%�,.�QPQ���#3��^�Z�����R2^W$���o�|AEIa¬�v>VEC�b1��q^]�Y$\;p����Oh]9]��m����6��f׸����e��8&u|��H�9ݛ���y'7�#UF1��Zb�P?���a�����=w�Azjs]�J�ͪ}�n��e�%:ZQV-����:ʜ�cQ$�a�]7٨f�X����!�ta�Gh��lfJ���;�cVf�{�.��
򱕯:N;�ִ��ǉ�`���Դ�J�AL�u�̄nkC2i��Hh�[w{��H� ��D<s���n�s���չ���w�ٿ�s�\F�ž|�`�@�q}4*6��k/̀ei#����!�K�0��`�h�v$%$6�>x���0�e�#˽nRB��^Ʒ��ȐI�"�i�8��@:w�e����\z�<ϻM�#�v�`��+�����ߡ\�s%�J�VT|^��Y���\YZZ�V����XU�\�qD��ɌW(5�Su�y��	��BC��|p��[>VC�x����N��:���:1QzH����Cޑ�bA)���ߗ�m���d�qN��#�:h�����=yi�#� *,b�qo�]�B���n�S���'�Ѕ������|J؆)C{�_Ft��� �8��ɺٹ��?w�9腾�a��`�%�Ӗ��o�Ҥ_�QW�ENW^��b�gPC�)t �i�~�H����x�X0rmm�#S��W�,�VP���@���S�"�,i�� �X��K�Q��8�n܈<�_G�.��l{��V��J�I���Ev����
��;m�o�x_)�\��B�e��_���3b���נ�Os4��?;{J_�r�!��N�7�_�X����j�D��;�T�rF3+#��*u�CHfj����eي0���y'�>j(��3���g(ՔG�x.����*QRTʑ�s����"�a��H���Z�(�-�G���lT��Z�wq-�U<�%���b�����/i�\ G��`�����>z7D�t�`%�E����w��O�}}�c@�j�?�ܗ��{�i�|g�'�UG�dRKT�{�+B̏�өl�B<��6����9��y������sǊ �k=�@�5�2C���b�d�����rٗ��)����S�퀌=�>NN���7�d0����/aAĝꩩ�rgL��(pg�;��%ќz}J7A����o��V�y+s�`��[��B���������Z��Q�J3�Y� KY���3_f�E~_k�N�uԄ��^�$�n�(��V1��8�� ,�2��bp�������w�y@��+J(�9�T2�gjb��ȩ�嚯���@�%z*V�}�H�q��C�HSP())�7�N�d8�
��}�@�b�T���P\(wgY'����Z}Lg����;���w|_�+������C�6;?�q�?j���P�q��[T�	���&Ȃ�Z][�<�U�C���;&��^a<uVP A�q� �u�;&��B���m�X!5ԹW���E�1��~�HGg��Gw	VL��~��Z���|^^�$�s�Wy�����`�)��e�^k�C��H�B@:�|G B�\���l��q:@�uj%�w�w�--e�3�:�\�1%�w�w��tO�2V�b�Nþ�'�b� -�g��x5�"�9`����*�z���tck��a��۲EZ����H�\~A�	�ls������L�� ��GHx���]RXDď4ekck[Q�x�laZ8::�h~)q��b�@��H=��� x&�,8�����1���$E<I;��S3MK����:5݌9��Z<���鮾����,.˓�<,�W>T�ih��7
	��V�s�_V6f�j�BxhCz�n�bj���h]���KNƒ���Fl���i[pmJ��p~M͜�EU==�
�)(�a��g 8�Z����"��EG-
���d�֘��N�
p�윜��ME�C�/F���2S����+���)��yצū�7�|����uH5�-��KIm�-��!�]����za}k��<��V1�S;��6��r��Ba|�.e���o߶U-fv8l�4K��</�_�P�) ����]���#d��hJJJ�H.hN+��ut|�uu-�V�E-��82u#l���jzzt�5<���M�Q��Y,��7l�or��XR����cu��ϊ��P�{�
 'LĿ�8A���VZ0By�t�j1����y��������ԗ؞h�'��{Z�B�O�W����"�ʥ��8:9��&�A�t'ڦ�_�VZT@;�&�O�S����q+q��3��Y&h�Bu�u��08`s�k=��e�^�ٿf$�r�!hU�7o����TVAlZ��⌄�	ق� ���jRqFd��)Q֘���������׬�uR��dJ�/X�"3�QI�Cn�6t"m
�H���� $��q�S�אs�R:�_hNPT�a��Q/9GV�)P��J����/����8�ֈ}�:iNCM�6�r�JM�{sT��m�v~~���	�):�}'�}VRS=F���F��A�$�Du)��HSs�8��� ���[�z������&�/��10gN. c�]�����1?"�)3K�(U^�Q@x$^K]%	K�KjF���H�8y��@���ylՙя�pE�CȎ�O�l��T#Yt!d�d�~|�7��4�R?:#�y��ǐ�,v���X�aY�Yǒخ�ޒ^{N(�1L�w/'�"�g�������"���o����I����ooo#����B'F� ~�UgQ���	{�"���,���vG�]���%�&f����RX�d7e�%/���i�Gδ
�O,���Ǩ�H�����>��6�V�a0�)P��L�˿X� .vgx�u�6ۜܟ���l�����?PK   ���XR�\"# � /   images/16f29068-8fa2-43fd-94bb-aa3b1aab738c.png�|eXU���B��Hl�"���H��Ҩ("ݢ4H7X` ()ݠ�ԢA�.�\�t�4��Xx��>��o���9<g;Y�9���1Ƙ��/+AJ|����J޽� �9����m{�\�y����-Iţ��zT�5����]5���&�0VT��ԶwTm,lt��1���6�u-��-����`0�0��o*:���l��b���/������q���<?J|��yV]"l�G��ׇ��?�8\���ʹ�>��N��p�+�{�+�=�������_�~����R�sK��0hb$��������!]�\��|1�����q���q�.I?�_�~�L𿯕�pZ��E��G���;f������!
�|���X|��`y�<"����F>�������j��Tv�q���FD�=t�{�\˸U-��k�V�NF+p��G�ڗ�+]�(Ǵ�=���}%��|�tB��I
~9O��K�\Nc�u�������}�������\O�D�[��oԖ�����
����}Hs�ş��r��8�\W�4�DUTT�$�ns�nľjܑ�����{��b�i�:0g?�cձ<V?f_�fr0C�U��q�+Q\�~;
�c�#"]�%�[��6�N5�]���^֥2��e�(�%�w����{:�{0��՟b��X�Jh���v���Tj:"�pn�G�=�`�?h����M5��AÇ�a��.�ka���i�_}����4�*���硗y�%�ڹ�m�e�T���S�99<�cS�0+̼Pre�Q��r�:�:��V��R��\�~�i�`�KE��Zƙ�t�^d�n<����9�﫩�����x��Z��?u���.q�J�<��O�C��~0����1���vk���I�q(Yih)`7ߑ���S��cf���{�/�n����Ɇ;� ŋ�������M[����ϲ��r�Vʨ�4b���9`x�G�>|8bʹ/�8·Vp�����T�]���G�]��VK����rT�:,������m�i�;t�(q^k}K��DZ�os��X#|���c�fL���YF�;�,�rg�DN�d���zz�	�����_t����?6����x���kf����^�r���oTЇ~Vj[^��&2X���������I��2��!JJ~��gW�v���v�3�Jì,���y��%�K�g�&)�����X�R�o��� H���)�@��E�E�8�~��HKZ���*萞�����l49�!��yRN(F-�`�Sfjj��{��=�U��|-?��ϼ���րo�.�m�|�1^��r�4kf������t��7�\�9~��)WY�j�(�l��1�����w����;�q �`�q9�Sz̤/.>~��u�FX@�w�QJ�$>t��7��".˄�ّ:��I���1�m_��.}s�QS[ے�_����.�U%��QO��7��#��.Z�~]�͐�Z��_�^*F�g�;��O2Z����UWDE-��֎���O��|�Jj��2��}[&�ʩ1?T�?�ՠ�E�}�'�\Ŕ�m���5J���4�6�xJJy��]��z���A߾��uPq:'�(��f{�Q����n�������j���&-(���w�{��VJR�YH\��CE'��q�#�%ڲ�>t�;V���4�c<<N~)�bґ�DLJ����Vo�M�̼O�U1͜y7Z�k�f����	��}5�{���t�>Œa1X��h�VQ������h"�`m�/��ā�yb������]���Q���8���V#.�Xz�Y�i�y�~�*�`��f>���B[9�(뇰��{A�M����P���gy\N��&I1���2�~�R�?Rv��.�λ�jZ��C8u����lK�E#�!������3���D��sɁ,*̬�h7����젦u���ʥ� ��?��a�����]�g�N2ʶ�l�����6�fp:�Q�:Uc02���p���j���"��������ǔ�n�|���v����o����s���+׮u/_p�o3�#Ͱ��D{O+�������^���]?�P�Lll��K���z���Z%��3a�	��&��v<�)x�"b�԰�-��*���%Ǭ�*�y&J<�z�6�������qj��sv�B����P^� ff��tB���122�7�A�]��=���t���k�`�3MCIK뉔��]��� 6 �f���KHH�̃�����X�S!�K����]{�UHZ���c�D�b���`��<�mH�0 m�֡b:���U���3�K�$������_�8Ե_��1�@�8D�V5''�ߙ�e
m1n�}�����ҧ�����w�+���9ߙ�xո�0�����ry����l�B}0Gp�T���P�t�~7:�����S�6mfҰ� A��c��������"��&���55S���'�"G�f��M;S�mms���0����Gp' ���g8{Rղ���o5G
�t0����?*�G��_8�fa��W�ڟ���B��`8���}������k$�Q�A������ܩ�$n<|���
l���3�R�K�.�@:a���%�F����n�9��75YZZJ/u�J6�,�PTS3�ō�����L���з�ii�l_*���Ƭy&��h�d���I����<�נ�jwo�[H�D8�;�~��K&JD�Ν;R���j�F.���x��F��s�>�N3+)*�j~o��x=L�Կ$�C�\]�殜\�m�������z�I�y���!�֗�0�س��^��@��F����
����]�2���܃��r=>Rq����̡�������C�=9�g���<h0,��j6�_���ryZh�T����l��H���jzw3)m0���cR�^�
�#�x���?(��c0^(9#�V�����P�&�������9����.�^|#dvk�G;|�����?,��r��K���$�X��͸��ı�i�~I�7n�3:3�]��~��[�áQ\�u�p�}O�|�ΝW�!qk3]a~�?~�<���#q��$�.<�D0�����T�繞�FK�*� +�|�J"��o�(�H=1DLIE�~�1��:�P�l��+�[��8p��T���h����G�W�3^4�#x��YS�Ы�����[k�%t��Al��iOVbi孟>�G�;�Ȏ�z�C��2���͉�.pv�����vS��s�.���Zmsl�.�g@e~���oQ#y�B��4��C;��D*�(�E���!$d�E�?IgBogci�5�]��鵑�V#U!AS�#��J�#�����J�ZԐ$m4A-�@A�-�X�k/�ˉ��<v2�q��� y=M��c� wp������DUs�F�O���NLL�wgϣ�o`U-�/y��{s�qz�}�%.�_v
E�7h�&s�B��J~���A׸c'/Or�oދ�nmmͱ�SG��4�^4�@Q�}Q8�z.E9���ʥ�i��:u���ԵI�>ϓ^��!Q*Ϙ���{e[��$/�w@� G����F�����J�'���(/�6T�>��75� ��S���M�BР��@RY����U��{io�B�ܽ`v�'���k&
�.��q�&У�"�&'ZA���
::s)��=��/�#�(�c�C%[�kE�mW	�����˒�~�/Z�����Pq�g�u=�A�>�1ϘXr���9MD�:�(*C��`?��xQ"H��cAAAVOC6U=W
�*C==����?�ܵ�K�ҹ��М���쑯}s`�߿�r(��@AW7Fܗ�9@,�(�X��1=��0����sXSpQ��G~��zi���Ʉ]����T�E��'PY]�N��(ϵ�u��mU-�˪en���h�`N#�����������˗5S��||�7o���K�X��ӣ�$�@aqw�S7\D�f�>Jd.3/��j���2����hJr���J�N��k,�%T�)i�]��~v�-T�ɏ�'��[ ?H��g��o������:M@M�|�y=!�J��x��T��3�Q6��p�۵��&�k���&�N`!��]�b'`=��)�(+H����}�������Yp��A���|E��;'	��
߆7.�m*�X�{[��[/ʞ?ޔ�-����"Ք�y/D�<U^=�_���.2�N�5��W������EK�s&!!���ᷯ_߿{�f�hr���&%%ErmrJ���|��5�>%6����>�y�s�PO?m��P4��/h�f&�]�n�p.^!��� H綡`����ի9P8Ǒ�;���E�jv�{`�L�Z��K*��J
�����m��.�C��l���R2J��n��<<���2�zd���:�(�>��#H@�q�ę�B�EWxxV�	�-9*ji=�������fm߶�JX|�С��{��xn�.e=��.�	7�q�Մ��qbe�����䅯$�r�p���jߙ��f6���4@���}�N�,�����*�������ՓѪvЭ�� HH���L�3��\�|꧑��ngj��AK �Sm�TUNc�ɀ̭�8_i�C�$b�(9:�T��Vյ�HW���յ��9�/rX0 O�H���yii�ظ89�-���� ]*��S�
�Et��r��NNuuu�;V��Н��T��:`K�D7��'�N��_af�����������$���i`Ev��}O��J��U���M�z�8�|�R+������?�`�Tmb����y���O��y"�P@���=���q�^kW����ȭ����Z{3-�!`l�� 6��0
���ϾH���Ť%�r��EZ���L��I�SK�G�~Q��P~i+�jq��<F��m�Ӓ���.���n}�����:k�w��K��h���9A$XYYY�@�üt� �� �7u�-e�f�V�	f|uVRR:�sS��$瀼i���YT�ǎ#�s�i~�F�Wto�E8�/aw�*åKW�����s>�̱�A*��`H���M5��iE�vV�˟��U]N�x��Kn���W�ѣ�_�~9>4?7^IHL��311��Xn#���Ҋ�e�!ۑ>�ټ�|U�"zs����&G|E;�sD3F:ޚ��Z�\�㷎�N�
s[/�2��nٖ��q/	b�HLMM=�t�%N"�3�� 
��7��W'!�E4��\��:-%`�vM��ׯu55�G䍍��ы�nť�6L��W#YO�8p*!>ŵ��i)��a��J)ʐ�/}IO�_U2!"����q5+�f���n&�4�@�l�����fuBt�g�Xd*̢����W�����~x�(x'�_��)�le{#�W,a�e"��P1�>q�i�E�i����C�~�CCC�����T�~ǯ׈�\�rWRRRJRR�����ve��<�����H ���ji���*q�m;����X8��营!36�磣z�������s�����an�9�5K�����,R��|�ʞ��3ok�@Ґ�6��Ӽo�@l���].�d�V��1�'Ca}��gD�_�m=�]��-v�����}Sg�p�։'��䂫GZ`�@�Eh�,o �i�	2�a���/O�/�I���*8S�_.���b֚��J�s,q�����?9�=S3fm������40@?��	�e'|K�}�w� q���OM#KF�[k[�)9�S�QBw�W��3>}Dp�j����g�������Af��T��?PP�(�3-�dOav�Խ""�����-�H�����6��������I����h@}+_D�1<5/����e����Z]N!�.�/0i�N��u��I��L��!|vQ�}o%��3��_�E	�I&`���=0�hɒ��"�"���M'={�ғw�~[	YPdd:�B�x�DC��F�ְ��Iroޓ��8�� /��
�
N��0�)@.��^	@����Ȕg:�:PW�z��>od�k't�i\G��:P⢤���N�"�֡�k7����Ғ���ƻ�#8�9װ��)r"��	��<��Q���y�J:�c6X�%�E&��t���+���,f�ܷ�܀^�W�h~�׊vMd�O�Ҧ�=�L�dg��r��TI\��^�����\�^HKރ#���k�#�5n�/��J2��[��K�(ݒ""��y�&�a�I�}{LG����ߚ����;��:ۓ-SK�z�h��)�w���t�Q�)��"{��\�rC��M��`��ЕJ����,���l칡|Mv��6��������߿����ݻ�����%�_YE>)<i�hru��@C���9���W�˗/�,,m*:O+_\>1F�)~��J�h��� z�1�����������R�r�zp�t��DS�Lmc]]+����f�'��H�YBJ6�JGA��W#k��gG6�	m�B��<;Ƽ~����w{}�[d�LG�C��\�]�������"�E��A��G��_?Uu��^�	���D�u���0�V��eJ(�� !�:[����0�G��o��QIЌ{h��vGǐ!L�D��m2����!�~,����R���[(?Em�t�ҍ[����a�::��g���YT�����'�?}�B��O�r���8{H��K{�:�ŋb [�ȶ�v�- p�����7Z	����ʆ�����;z�;e� ��"��{r�Y�j=-���rZ�w��	II)`���h����%'WY��u$ܣ���7�J�T�J9!�g�9Xb#[es�t���d����A�<��FO��U Q{�4�_��^�[}��}7aL�c*O�\��w�w����8IFV��W�жA��m=�˔�o^=��G�>;,��6�wJ���FC��c�@�6קyRY|�!:�
��/�{���X��l>���Gx��X"E������Q�+.6r(q~�L�Yf���55����s�l
Kz�-�W����E�Cq0���$b`�P�=���!ܚ�<��1C��g���8p�Z� ���@�[��2�o߽k+vZ�����߰
�fҖ(���=61�"�%�Z�Ձ���qE,h�Zj�$jz��(�t��n���lR\�"�'�����klT���-X&�I�����77gg�OAye5�<����t��%�kW����͏អ���T�~�V�|�x��a� �Z?G�|mH-��&)P�~E�vvs�J`�U��>����!��"ӡ�g���B�C�]]������R��/����vR-�v�y�,��7ڀɰY��G�5q�='%-̓�\�!� "l��SV��9JL�@Y���C8����?gx�>x�P?~<Sz7J�=���LD�1F�>�R���2h�|"u����,��2�A�SϷ�aB�����������CY3/���6��`�@FG������'���9�C������XQII_j t%�GI;~a �rJ��d033K�N�a3�mld�����IMe}O+�=�;�p	�- ��7ys/1"�6f�E�g?���׺T&��\qo�P5�K�~LK�� $��en%Lj��d�qQ����hT�jd4|�,ʟ����5j�����	�o�,מk���Mf0����K\�2�8�%��Y�AvO@H�`du<uU���Tp%�k �"�~�]&@��z`+���x�J<�L�(��Bq!O���Wh�`v��@F6� ��P��v ����㜖^��e[�.��xz"8s��OU����s��
�~R��:�ߜdL�̞���삁U�ˀ�09�y��x�kp���e�Iz6�Ǐ�0
�A��^)0��ǎ}-$c�QN��x����#���� ����HA��=�B@x�_ݴ �J98D�f��p�L�Y�'>q�m��HTw��Nh+��ŋ2����������ڧ��!��X1��lmk�5i��'D�yd~�,X?����
��zv���&[��h�z��Qqy`~�+��5d=�Y�$Y�ǟ�Y(�Yt�? ��V~��O��g�ނ������s�v��H��)�9y��я����V�d;ʻ�A`�FO�x_���P�7w���7����I��
�������dK��������>�w2꫷!��3C�!�{��&׳y��;t��a#gh���d��� �T�
T�Ϋ���Vd���U�v�`��M���8�Oc�e�0���9F��H��~���p�|���_$ �cN\�t��u�MT��_,8\fa�"�h�3�M�)�= ��[��`RC�����,����FJ0�M���壶q����6�4�8:�[[[�c-t�e}��ҫ٪@sz��ؒ����k�«Sm�`�ύ����>�^f�u���{������J��q�0��������ߪ���I���f����G�y�=�iU V�uݰ�{phO��ޠn�P�;米�����ʨ����%U�+a��
jHk~:UI���P�I¦]��\���>H3�Q���-�G���k^��4�zpR�l���,��ϿM�C�j_˾G������1�e7�ͥ��^8yA�}w��2v���1��B�j�x��� �n�2W���`���	��w3���G�C@@r�h�l�2��<�_P�X��qo�#�5����-�b��	�Ǐ�-9Jמu+.��z��|Q�S���Dә�z�(��l:��e`8�H�_aJ��� �YX���͛dBBj���-J7�=�ՓR���G�gB3VZ$���7^��F�"Ga�O�ѥ���l?|��q����	>�=6:��14����g����X�Jݰ���Fý��oN&��eT���"���<����T��^������P�% <�o}}�2u+�!g�%X��L�Q˭
OR��%L��D���/ᖡ� ���Ǿ!A�!��]��.&����8C��"h� 4��K5ݛ����oy�ud�"L��&��b<XZ�I�(�3n���L��)z~ j��4�$�c0 53��M3���P���������P�:uJ��E���ϟ᳌S	w٠8`�g�Duc�jZD�����̱)@݅�޲��N'ğ!�.qFҜճ1C���B�
E��`���7翼��\��_���~y�?c���[��#G�(����$�RS3mI���@7�`^ �������t)��̯�g��_�-pJ�����b%�~�C�A;H�v�1��<<ɾ�t*��0c�],Im�v�c�Ev�C���rssMMM�oȿ��B�p�g��F�����N��� ;²� ��o�+\��w�_�4���?���3���}���w��%v������ٷ8��t,W��4-������ū������L}��(L�}�w�O�kega/�����Yq��DD�8�IFY$=(-*�HB�+ڡtH��.wP����hjbR73=-���A���I�%%EPQE�� "��Okjɱ�S�u���G�����P��mY�y���R��'�S�ґÇ+���>EGG���8AGC3k]��}N����}0�(�;̍Am\E�Ӏχ�?{�'��Wr����2]jz����Bv\a�V����df.ܶ��v���������>n�ޅѫ�e`�61_3}���ZhP�X+:�U����{��x��4�9,S�i��%�}�E��?�:9���#{w��m���w�h]b$~/�1hdmaP%2�cG͹�]�����W���K���FQǔ�[��ڴ�;��t��0n�^���q��X������?�����ѝ���F�o U�\��@#�L�.��M2��ȼ��sn�z���+ܱI]}�o8�Ӕ��P_��n�0����qs�%;��c~מ�[y��c��d�i��\�Jܾ�s��uw�}}l_H�\�d�t�Ѓ�'��W9C;��f����3���le��L2�,� ��;���ԧ�D�C�Â��2�x���w;2��d�[{��,F�����;���ܼ�yw�nTέ4�,`5!�^��Spp������)�� �B�t�@14�Mӡ�!H������-$s;D���b��ݷ:`�������,�F��m����{��X�^���� v�Xv���w�ky�穋�R))*��,��� ?J�4p7_ad���3�U���o�B���M��Oה�� ۽o�+��V�(vٷ��-A��_##e��^�Tժ� (����>IKN�R���������!Ӡ1�_���ST�c-���?΃�c�*Y����\Ft���c�o�!F�*�#.]�G:	�тদ��. ����6��(���n��1����wo��n�����%&%������z�U����ӮÔ�� l�
����A�cA�����stt���Y7g����b��cs���Q���֡��w��W8j�޲�.x�2�l��ژx��eMII��ty�+)��<������� ����uzxj�ӥJ�(�.�W�������v{�7���F�a�E&�"B���,%�_�~}"���/��8�mf�u�{:�ï���/��d�)����)����/�����w����Ą\�5��Էo��A\tq,X�4�39����������J��X<�V�Б�=W���PX�Aו��n�τ��Lw���ef�
��ʆ�Ye�T�-//��φzROqqz���!l���P�7�ͱ\���<�~���|��MZ���Z�I��U�ߙMK� ��7�tf9�D�PQQ��F�y5���5p�7�e	L���VŬ;s�F҆�1���D�6����J}@�%�(?2^΋�vjXpрN&�f��݁?6���3G;��j����
ZA	f�:1f]�������o5:v�����Ԕ��5;�����Ҡ����o��ٜB��+W�|�$�u���/e�U�%z��������uy�  @V�C��C�!�:���"���>���-JM5���LS�P��\����olYZ�j|<���%:�VH)���~ѿq�m���U%�>��4��9�W9
�۳�Y=g�y�>q9�4^_�FD����\�͛ϴ��.����P���r_c%'	Z�CסTY="/))9�4R}�p��>@�h�+c?)������q0����4���5ݻ�����*b�v�,��٪�ie.�B��+�3�vA�.�9.�S,c����z�������傘�1�߼ys�R�����������8w���K@k��>��������*[�0�)z�t�Dlssen(S�[�f(��q���L�H�'�jZ�Ipo?!��"�Uo��E.JĤ//:������z��T���#͑.��~wC��S�+KY]]=!..nm��|WN.g޵�P�\��E��r	�ݭ7Ër`��f���j4��[]̸͓�`Q����(�/p钞��٬p({J��٤�/h�me�Q�q1/u�`Ӌ��r��Z�jkkѱ� v-t��K!����&ehR\���
t�g]φ?�)S~�b�4��rɰ�9���փ��s
�Ωc�q����/����S*���u�ʕ׏q�bK�l֚>��7M�y&(ݕ�D�3C����	���6������;3t���pD�=�,D�:SH��������ѣG���v�<NL�
ڋ�Uh�,���KIY9��iWz 5�t�#�-;�|Ok��?��>��(�r/>op\B��?{�<��{��0�в������}%-��]�v3o��_, v�l�	���p������|y��]Ni9�z�??�hҕ��I�j�N@pp��놯��>7�(ZU���L?�G�#��m�f��A-]����N�`Q�3H�=�:��;�4��>8f����99��^���,���� ߃a�P�N@(j6\��8IC�V�t������e�6�fZd�	P0x��$o��'mT`����\���GF!캅2ڔ�;D,aV�cll����ԗ��E$3�E�G�^����D���TR0?+3�>[����[��פ�0[�͘yO�����'իX'��חB�ļl�^!�2/���]��O��δɉ�am�Z/U͕��
�X蟮�t�����S�/����3����qp�FP�����z�c]``^~ND���@~IIA�[^��P���� Ad��5�k<]����,��)@}��z��	����10e�9Œ���� &���/ {ĝ��X&'�� ڍrv�DO����nՔ�t�����;��� ����g��l�p��ú��j�.@���DS���0�I/ "�����1����ƺ(ZI���mc8~h7���A���!�"��r�����&�����y��H��b��V���L�^��5���.1�l*^�E�7��NC��z{����������uttD�ʲ�3������+;<w�f޿�@���
�d:�!8���F:��'z�������瑂(���@�S%���*زO�C/ȫ�u�����7���-x�;(�⪙!��|O+b0?�@�߾{'S+u�^>�7W6F|g@ yX��e�y*���g�(~����U�VR�0�ֶ�DS�\��r���k�dŭ ���J����3���JBCϤ��%��tN�%ɕ���P�WVW��{@��-|�E�KA�6Ʌo���a�C�Б���� W�����y��}YY(>�B������ֶ��ly{��-�1%����e��EkP�鎔`<�tI*�/�t�WfTc��e!n�@Nf�n.G�wөFB�pD9O��Z���Y�n����1��=I�v洶xD�o���c�
-%� �v�����p$~�<ɕ�]. >n��@����$ڞQQS������-��M�ݓ�����G���G�/|~m�dY�Ul'�%m/�3��P����g�^����e��������A�p��Z���fҷ~K\�[��t)Qi����1Y�Jq�!\��jjЋ\��j=��R�ٹО���,����t�^��O��S�G��	7�=�e/ѝo�knk):� B���<��ě�������;ZZ�a(�mp��;;;���MZ	D"���Z�911Q�H��G�T�u�8����$kZ~;�%eR���C�<�w� ��U���C+��+�I��6����}��'%9�W������#�^�|�$	��r�'$T~�E�b�n���g9�B��1k�Κ��@gy�ؠ��"��������^��4l7��OL���W,"��J]7?�7����-�&|�q�nZq�;��CЙADD�	��ݻ?e��{�^�g{l:��M�v����/���SNU�z2X�4j��h�$~tt�uI
�>g0�Y�cR�Esy}� �gڟy���\%�C����;2�@ȱaBNY�ߏ�R֍,���ݻ�A���ж=�"��\`Ɣ���� �M������Q�m�/a�U!�6D
k<x� G�w��+p�o��뛛�U��:�,���ղ�&�);�D�7ߠ�8n���(�'G r�d�����u�2XpV���������f�^g�Z�=o
��g���(�	}D���*�9o��į��͑��]i�,<<�7wM��P.|B��0���Z�i�7�A��EcQ��z���z�/�"�TR�xAD��{���P�������޳�w�^�I�q7�	B3T�_9��W���#U���`��*�?[�Q�B��H�L�󭬷�g��6
ϋy�@���:+R�3�iݦ���d��;e�^�LCVMY��龿'!( p�s��Y
�"��^&�W05�Smǯ�������<�|{2\�0͞<�q�6(M�믗������m��GO2�z�k\�|���R�kJ���^4���L�6�_nm9�噅���nT��%R��m��_�_(^�t횲`��[翤��+��V[�v�?[gg��hN����*���� U�o޼�&� p����1g2���� ����j�C�+�����x�1��~��붒�����6_>�ݮ ���:V��M �,�	Y�NH^�o�9s��LЀڢ�R�uyy�G�>��� {�� 2�~�����B@/!��Ͳ}�N�����C:l����?e_T�f�}�őڂ�H� Бg��њ�Wmƥ���4Rv���Z�7{��sB�d��5�u����0����$QDz3�ٗ.^�T��:U�c�����f���|��[��?/Vc��;���*W��\�5hǫF��-�x9۰9hu�v.�������1�Yp�`f�S`�r�F�t�d�w����4������n��<F@eY���{�nD2���P=:66f�=wut|\DM]��y�Xr�����z�`º<�OS"r� ҳר�J�X�`�7�rVNS��v�����q���ύx��v}�^�ݺ��#�޾=��Y�����#st/�wƯ�"��� �EDD����㱟U埊���f�%pp���4
�6�U�ް��EF÷���,�_�d���T\\�{/��V������\�-�G�bB�%�I
a0KF,��=S��Yщ"���LvE������l�N��}�D���?�����ã#Z2�᫾�N�����)��20o?�e}^���T��mwj�_.��q���ꙓ^↑N�$���q�<<<9� ��EQ��sYiZE��@�M���L������LI��T������x��w�@�́�RC4�x5��-1d��c�pc?M��5���0Ғp!=��A!���|��OMc#��E�����nO��..//���5\R�h࿿��pm��z�p~#�e=:�ʽ%�H�(��������a����Eyyy�ʐr�ED��m����)���e����[�VUpr*H��6e����)�p�>G����G����0��>�]澟fڙZPg�%�u�����iPL;�:kR����X�Ms `a�ԽG���\Gs�dۚ&)�ݸFtE%U�ꖮ�n�=���lR�}O��H���#+���jٗ����� �����!���m,�l'�߲�kn�b:��	�1L4ci�1?��`��TH�Q�|��X�~pŰj�as������\����C���\n�7��~W�f2]��ZZN���C4ő��ݠ��!�]��\�LA��5�h���z� ��+ͱ��)	��_Y;L����8wL��[����VɫBb��0����2��v�WR��~�ldkn>/;wz��ԩS����:�_��E�q��U����r�M��az�Q����4��$+-%|h�����-�ZE�_�PPR�K���xٿk�י��K�^6�D� n�3���+��c&���� ����p�Ϋp�@�`hjH���ѻVVK[^�﫪v'�mg:�d��V�����b����L���WW�*K��;3�9�s$JJJ��ܦm�2�N��߃ۦ\�@0��R��7D#�>�X�#�O��c����ģ�>��8��w���E F ���)�O�5�@k_����{P�V�r-�//߂�)�Lc�� �x*��*S q�N-�D�ů_��2}�ԛ���}$b �Lll��YY���9�8�����0-II�����`T� |��?��F[$�)��;����8&"]����Ҧk���cG^x�:�'�R�h�"�xT���r����VVV������0���<DW��N_L���1N�H�Х&ɗ�"ă��ٕ�����PbP��q���������Jl����J���j����:�N����L[���{WJ����YiN��.�\a��,��`$����/00!B�sU��Ý;��^K���-s������%��&N\m#箛��=�mkJ7�]����`����}ѹ��w���;��[���$Q&,񀧦Z~Y���vg�.�����!�OȻ���U��-1�	Y٠��O�l�/�LDL���z%-��aK��!*���.���G�9W+�a�y��^��j���
ڧҸ�~���ى2Kw�]4�5%$_��+�IT�?N��a��Ĳ���-Cv>�7 x�ȿ#��(�e�r�k���0�.HӺ�Q�G�L���ₕ�^���6�'i�$^��~2 ��%4�ŜK�յ8ܮS￥������i���96?X�^1\�fN��u|��bt��J��N��k_�.Yh����dN+��I���k3��X�?��)ם�j���xA.r����0�j��:���#������t�Y<�>�I�:9x���fQ���ߏ1~:C8��E��~/��f�-��6�ϸC$/A�'�X���020��=��`n���W���$؂���珐�[�9�������M�/�
=B��ڂ$&���S0ؔ���$h?������y��m.?44����8�(-��\n�w0��rj^� {����ز����b�r4<��L`��":_�hܣ�K#�^�N�0o�:D����h�̻���	��vqw����Z�R���1|�h�&��#F�k �nV��k7'8�g� -)�
D����[?���j���?�|��\N[7ɰ}�S"2�Oc�FX�@f
ػ�g��w�Ɇ�V�?~�02����{V�=_�����H�l��O�_\� \-�Z~MB'ԍ�e�sY&3{)v��R�:�\A)�j>��3��1��<�`t�;BW
5�MNT���5�C@R��O�r��2��� ~����P���8B�^�GM{��7��b�uMMA�(��?�h6<��\�v&K�ٹ�U5���s�MNO�U��0Ud@��)*Q8�+��������8�n����]�
ۍv������Y�ٹ�>�]3�ʊ���N+��wM}�zۼk�U������U�nN|B9��˛e��\�&�>:1Q�o5B�q�|��߿�ҫ���Spgels"*x�Wt �� �yy|�F?�w���67�Y�Z�1�`�����ҿ|aR��7���§�6�r�[?��<+E1Q͔����ׯ���}1(v���s+l��&��7Bb/Y���8G:���$H��*�QA �6�:h�Q���Z��DG��@�<��&l0��Nˣ��f_!_�M4E�`	u>���Z��,���v��I��N�XC��j&^���������c�s�#U��:�	�ppX��r>󰯓�`����Zp��dt�v�.---��׀���+8�G�}E��f��mms��gҲ��.���]E�h8�ϯ�W�vS�����>�n�f�II�Ů���"��[vW�Ο�)X�Ce�A�ߪ�ؐ&Z�$��q��k���	>EI�A����cQ8X.���d���k�7v7
�<�A����:r�Z��Rm�TUݍB�[?��i�r�����n�΄l�DBii���p�?�P��0g
$�k��v`��4�ƌ~TW�3%Y�yrpэ�]Y�s��)bI�`Mq�To��k�����≍��,��-9���S��ILJ���D�Cy���w*�Nw�_��蒑���n�[�#����K�m�m_%o)���Cf�s����g��={{{���l9�kkj~6q>�_���m�!�� #�đ9�r)�qwj1G�h�țVPY����^���k�9eTsR��^�咯���,�4	jL
���g+E�ϋ��'�i|�ar��
J```�k��{:O����;šJ��HH���H=y�䎸xUA/����J���АE=R����g�YV#�sX%Z>So�,��`B���U`�r۷DP�@)����b ea'�	͞�g/����ROSY�?FS~�<�j�ǋ��`��(�h`X�YYg-4�4�Յzٞ�]��u?�������Z������ 6Ts�#~BҎ^��k��`)
�d���-��S������w �܊ �D0�cxћ����~�«�;�F
����ͅ���#�frg��`�.��h����	�W�)�8kr�����Y�"��S�tŴ�e}}}���F�h����l�{��(�U%k�,鐫w�(�u����ga������@2u�%
���9#'g�|��G�5��>�H5���s��z��-����}�F(���K<�@3���V,��廇�|)����Eq��!�c3�^�	F+J�"h3҆�&,W���%_PPp�E��d���eIu�Ѓ	@R쁼|L�W���Uq�e}U����l�������O���Eh�"<�V✋--����� ,���#�'�:'��-�zyz[#4F��7��jj�3!k��q�w��t��ud�Q�%�Σ����,��mfh�ze���L�bL�u�H�x�`޽{�&{��H�o�iF��|�d��t��b�F�0�����7��կ��\i&?��ٴϟ����y��64�ǉC�ހن��u��r�\?� ���sk�j��|��*���U�鉋�F0�?��hn��|ę��-z���(W��������8���ۨ��
�xD�k��r�5��bI���p�VD��t��>�7��لp6u�󔭶���g���  ,?g(��5��k�9W��t���5 ��.�����h\��D]v�YIɕ�s#�x�Yo��۲z����㓓���"� ��?"�eO�Y}�t]��խ��[�P�n�C/S����ٰ���?ޜ�0��5��_l}w<�o�����Rf
ɦ����2����ݱGˈ�dš���ǱJȖ������s�_������s��u}���~_�W�C��T�����r����w@]]���jǫ��'�P�^�zU��RSmՈ`�����]5���bb����?:�{���:Q)�]x�ߤ`ύ'�ѷ��E����{���MQ��-3��R�˅h����ʚ�S�#��E{�|o##����*��	�j{LL�����/��8z��lYf�i�ؗ�LĖۉl&zzCu�����9�k��PE�3�ˏ�ě�����1�7�J�D�'���P1���Zr���q3K�_�l3{#ZL��5�#�U�7����p�I��P��s1��n�����r4&�`QҞ����}���J5�!�-:�2�8N���;Q������ډ���iz�@��;b�ѷ��ĵ�p �;�bK�VrV,s��RZ��\�2�&I���=�t3�R}�yu81�P�U��1a7���=KbA�����q�d"����!�Oğ'�Q����N�M)^�ǹ�����\�ݺ	~��l���2M������`�5���ϯ8==}�̙���0������,�R��8��ɑR��E�i����ɶq�퟇PU!�t�`0<\%|��f��뭷��/����Rn7PM}�L��$y4��~��8?�����)��Ӄ�QW	�<��~�q���F�Ѭ�Q��h�0?�1��G�;���������e�v6ܷ?9W���
�<M��D�x|\�[7
g�E9�'8e�AѻTg3��΋+�s]Wq-�s���_|̷�'5�o���4.�@�%܅�oWёE ��o��y��ُq�BS��zz187� .� �xt�fg��ɱy��n].K�ZU�3�0h�l�܂����{!��۶@�����v/~B�G$|��莓Ԓ�,O]��T��'�� UUU5	�(�Ք�ɿi�[USs�����~a4�ald��Y&mk����H�A�D/��� ΀�{�w���FG�#��j#�C{��]EE=��t�9�S|�?�T�`�d$%��\c��/�%K���g����jH�s���T��ʿ<�c
��o��<	J��#g�'1L���Ǘ@R<�+��ۣ�:�vR�.���9;0��Q�dPL�@������'CCOݹ݊���,7E�̓ 
�	�t�/��';���U�
�\+m����1��� 0�[I�^Vf�mtB��Q���fI���x\fp^�hҕ-�-�̣q��a��}	����ܾ$$�gt��B�+���}�~��&IjK��O���]DV��e+���T����|����R��V��dh����
@���̢�TU��Y�N�?��M�"v����.7�1�;ުNX��	�z�u���vh��MKX��zb��T�ѻyꝧܴ���0@�Im��������@s;O�@Yw˅	8�B��5-#H>�N���(=~�d��x�
7Z��Rq���W��ޓ�d��I�
�L�����6�ZZ��J����ж�i(�Ҳ�޸*׼�����`ͷ���3�Zl/��sa0}��':�����|�����<T'����Ƅ�H�fg�M�U��/�s�u�v�\��/%a2�h�wo!,U���K�����N�����d6^��Y����="�hQ�81))�u����Z�J+F�e��D��R��z[5C�b�q�	�ޔ�y�1P���4���V�<����j�gPFg�)�C��~12���w���g��`�ǡ@�-^�o<�Q���`��-Ӟ*�ڳ3:;{��߼���y%%��Ô�#��������y`)�9989�6��Ov��><<<�������6������7��&�ѣY�h9�յ3���-O�4CZS35l�9�~Ag{Z����ל/�t�*0�nDfA�Ɇ�\�k(Z(��D���%���
`��:@of�m��iiw��
�y�@���A�h��|J��(C /������.ްis��)��6��j�`���l�2 ��>��S��Y��	�O���Op�3%_����3ȃ6x��Š4Ի6ic����)��0cׂ"��H���|��H��6�ѕ��vsZ.o~��O�J�,&U̐��$76>��쥤 ��.0p�ΏB��9Z�,��
s,�_J^>h�nk��X�R�>J��v5kml�����"�Z�Kx�����V���{���U/x(�Z(H)�L���/g�)�V�9����}0rc5 �V����+�qÇ���vӕ��u�$KܸQ�զ�bI��W|:~�<��b���L��!��
��kK1��w�^4���e���2 F�[|�ٱ'�F�"�+f���8d)J�궑�Af��u��d(p2O���{�r,X��Ҍ+�,D�r������gYXn���?S��s�q%5���)A��4Mb.A�'~���l�aܬ���c�8"Q�G))��P�x�n����?����<~��h�͵(-������a'^���.RAW� ��0|�/o<���$��e��1Y�0YM��v�4��t �������j��G���X111�n7�����bH�%���m�`a��b��Z-��ZZZV��#' N4@i��s�$_���w/�Z:zv�R�<��;)����h����;m�in~�[>X���)�"Opz:ߦ���T��0�')""B1���o�+��@��,,,�q=�==���UQ9/�!��tt����䦿�f�l�%�P?F����`h8���μ���!tFP݆�����ÊI$��~�B��ь_�E�FW�.�����ՕcƐ��R�*O~���W����� �,>��Bk���	YX̬w�P>5����
D���Zե&af��GV���!5+kN)���`^�6�B����lkd�AL� �X"�4��3��6`T0��S
�Z��"�j�����>��ǈ'�k����̪�����]]eS2�̬����=Ӷ�;��m~��'�O�а{zzn���<zt����������k�U�vN.���b�����?~��=�V�����:cRvvK�4�g�+�B� T���%oc}e�����-{�"x2��Pc�3�\�鑥�6�������8�[�4dQ��y}P������y NG�xzy�|�rÙ�-��n��M#X�:�a�&I7�-"��)>�i{m�
��Ž�s��v�X���G{t���cbc��_2F�F,2����$����:��hY/��ˬ��{�yfb���kc�EY��z!|]q��6�Ho:��=RP��|�NLf�]��yj���_Y���T�dF��G�"�&\j�ꊮb� ~�b��d\aDK��8ղ�d��z.UA���=�A?�^��!�_&�Ro���UCc����w�2op���W���6���`��ƌ���hP�_2	��N����-[�+�ٽ1�G{!����B2��~H�܁6פ��}����F��F���� }Y��k���������I2�_՚��Ϡs�EǄfC�H�.]ZS �L5��i����N��΃y~�Լ^ohd�(�μ��8Z`��q��hk{�oS���蛗.^T'�k�t���ǃ�_B	 7@��XH�b3����
wq�!|
��w�]tl�zʆʓ\Qjʪ��ム��s�0�����-�6.OT�'�F�<Zܺ���FRe���t�ƫD�6��Q8�]�s���`O�7G.�D�����**(����Ԡ��h?�]+~XB|��W�+@>�^�zE�>�������ղ�hj���6jsԔԙT��+!��`��Zk),�斖J9A�9�	�!�g<ԁ/���j_�ٳh~PޓZNN�roSU�n�	8`��}sN�u�$���9/ ����a����S�~����e~��'O�@1}
\E��:��u�0�xv�ӧO?�\�<�q
�S36NЋHL�e! ����O�"1P���5x���l��a���C�
�.�%�h�ϛ�ƻy�ƈ]t�iOAa���	^,�#�����Pd9�F��d�sƸ	jpMs�VJY�w���w\&�D����܊C�Cf����i8��	1W=������J��2!*(ǩS�6���Ѯta[&��{�<z!�p}$�f�2�u2	���]-�d�Q�BM��ty���ƞ�d�Q�IG�tSm��/�uh����{���B�F�Rd;�D��g4��Cq����ۯ�~�زH=1]��܁̣���W*�d*��6�@�2��B��W?�ĔE**��Kwf���{JJF�� ����S�T�lޤ�H���a����2�3�ˌi�̯`�M.^�T���a�	�8R܋F���T~��ſ|�Eq�`gI��ϯ��w屩WlTV��SO�B�
�Ɔ�y	���۷����Q�`�\��(c�:>t� 3G2����nNt{���g�p>���ie��R��ٔ�����C�~hKRV[U\��W�w����ԲM~ʧ�����;p��)Q��+!6�>|K-��$�4���p�C��{E�����ԧ�+����A��3:��������	[)��@��q���C`!��JH�2���J��ϫ嘶��xC��o*(F@Wt
5ut�!�eJ@\8�
�I�Mic�#d|�e��
������1���jNj9�AW0"jo�B'~�o ��ε �+)+/���1�����JC�W�յ���ڡ�[��A sM��94Y��BT���{��;�'z
�@klN&�NCE3�S�����[R�- VjG�	<%�e*�4x0�s|�?��5Y�f� �&(%��[���mX_TŤ>���E;��~�����(B{����;R�rccc���+��s�q��\��˲ 6o3���h::��8���������F ]\y~��M��:;��]��~����a�f�	4��@t��<��]i���fV�ښ�U_��8�7�%�$ ����ٕ+�SC��M�6��~�C�
Z+o�5_:aK�@d�5���(n���J�; &��(D{fMgn��'??�	@Hoz�M�ҳ��Pu�`/�K����A�Z�,� ���V�K��ŉ��^߷W�?~� �Ҿw�t���y���1_�Hc+�4S84�w�<iApr�S|�-��Hi9�78�b�A�)��2(lh����S��П�U�?;;��}+t<�"���
6��&����znn�;⛑��՜�"��3��b\�ZڴOR�w�����94b�%2�O��T1��H�yR�����P{�;���Tm6;0��ou{� 8��B���ء����ϟ��\z���72ϓ"���e+�E����/z�E�S��Dݼ��X���K+游D��-��B���@{�{w�"ǹ��6fm�[�ܡ	imD�x	��\�$d;/�[�7o��̇^t�`��X}�b�W:T���&#�D5677���\Ϋ�����lӰ�ɡ��Na����ϋo,����w"�b0L7�/�6\�l��|F�;Ӫm�F�^P�~d4��<�t^�/��.�����y�;����� ��?���dd�t��z�8��/��"eL�vv�G�M����a.4���8��K�:{��h�2�E��a�y�8�OE`�d�C:�rP_ܠS��i�p���x�����t��DD˼N�0�v����`�����@\J������Kˣ�8�ص�y�	���Jw$������Q`��L@;�YT�Q�nV�S<���\BZ�A�5�����	Hױ}��J�.�v9Z��h�؝���eq$�"�M�4Z���H�C
����`��$1}e��YYYfO��Y��d����[�~"����70)�K��-��N9�-ii�X���[��V��*FR־3�P���c��8�0�8hҤa
2� ��vW�0it�Z�����b�P������l�����ݝI�����Fe�v��|4�{+�0�c�^���C�^���̌�`>!������b�!���=���eB��ݻ�#���M:��}i�<C����f����+��P3s�����)�oK��\���_�/.&�¿�OP��o�<y���8S���N��zS]���j}���ҹG[��MC$)�?�.Zm�-�5�~c�W��-��U6��ɓ���7���b��P�Z����;���F*廎��O:3Go@Ē��[m�W,E��:k�|��1b�W���B�E�f��^Nw�p^��]gA���4�oA�������Jܒ�?A�0?�e�&�������������n���̌��늁�h���˨����������� �9
�@ȼG!�$$�mR�G�~����H+ �<����+j�U�,��
�A*���׃y#��:S���M	$�[rr-�5( �6��8��HMʾ�x���`?�AG�43��l����T����[�0K��Uү}�wsske��er�!��n�zT~�����&MB�p����}	�Y�.��`٤e������TyII��4�|���gɇ��dx�L�?�����e�I_u�P���3O�>ʭqi�|�s��'�~�Z�2���z'�,C5ndfV�;2���ۛrs�N�enػZ� �1��tim]��j��E���o$�$˴�[���Q�^=d_a�c��Z� �	�VEi�bKP������S�F�F�eځ������ƚUTTcs���.7`��u�v������'(((.���۾��d�_�w���$5�b>�}��gGr��F{���(2�0�ٛ�@[��_�^:\&�0��P�g>���iI��f���]	�ޠ)�jttt��t*�m0M�͙�S����F�mi�U*�4:Yr�hdb�(t.`!�&? $�<:���^f��___d��Y��t� ��;q����M�L 4��'۪���I@��b�f���60��X?����Dl8�$��L�&��uP.���@o�<x�Gl����l[���(������<w|fzz�7d.�ilh����už��R��Y���u�������ŗ�#��[���G�"����۠�X�(c�Ƃ���r�?���I�D��(���h �������������P�V�I0�SjS��jhf�r�/|QPP<�?C��f$� �D���0�*&���>))��H�ڝnۋk*�ќD7�s��K�M �j��N��$m͝�X �eo�t����R��d]������ǿ~�3��nf����{��h�9�4��.�ۤ�S��w%�/�����M���MB�[���u��񺴭����pA�� Gh3Cggg�
ZW|᷂.z���!��?EBJ�X�i�J���˄3�ݤ����m��-.���S�,"b_�;u��,,�
�/�����Q�X�"�W��qe�
���l�8�u0̑#[s�\ڷ˒::�k�M=
	ğt����r�.]��HGhYs>p5&��� <~�y��^�2fN����mi����3�k-X���������hi^P��(���Ԑ���M	A� ����n��ډZ�@*Z����#�`�WK�^0��̸��63r�s�6��kK3;!��Eu0������9d�x��T��l��û���C����hi�@l�ˈ4��L7���&$o����ɟ�����4 z��� yk���8������Q�D��
�j�����r�ᇯ��Ê��4��@�N��J�|����F�prr� �iYYY��]WN4���R���ԏ
R�b�f�?C�>"kd�r�O��Bz5R��A�*S�5�CrK��/mi����W��:��x	�'��ހ@�}`���#�����ؾ'h�Κ)��i߄Oni��;ԩ��r�t��3t�n�J��h^[&��T�y:��d�ӧO�'��d��b5�Q�~����yJc��o���إ̬,�dbC T�M�Ep��5Y��%��UT�a��?A��vnm�C>T��ߊe�ֆ�ñ��I�$Xmmn��(���J������J���Zi��~d��W�@��JB��޳s=��5<��N����� �S�Vd(����}��ɜ)��[`�K�4��b���ğ�3�Tf�d\G�<�� Q*�m�N��[�nQ��%������==�*`��h�BMM-<P�ܳvR�d�P�FƁ�7]�""X���KX��r��֖��v�����C=H��$���r>q�p~�,�J�?Ґ�V���.jho{��_he�y�ٴl|�|x<#Ҧ�5d2ϊ_L�@�;ƾ���"ߚ!�h��3���u��߂$"��tV�����@�a(Hϐ�_r�j*��
���Cp��V����ȳ�0p�9��q==��p�1�{_]�X�Ǜ�2�_n����+���l{��9�m�	�P:�oE����YɃ�_U |`�:L�̪֘7�����c$r>}�-���up��k�r ���c]5�D�>> QQQe���摏�w/nv&d��:#�a��;F@��O�^N,�]YZ���e�z��$y����ܱ}N_����M1d���[��A}��Y��@���V0K��H/7�d11�����������C�,�������̐u��$�eR����ʲ������4��m���ў���m�I@�:���:�@
2�P�LKK�Y�T�4I�Ίz�f����W�[O[08:\�5�'[����B�Н'�I0��v%�e�+�:��Ob�322��_�!t}����u��FU�ƻ�A���l0���/�I�^j��{ޡX��¨��.��b��֬_���Ɖ�S=�`�x�:���\w�����Z�+V�&~�b(�C�<E�U*�+�~��>"q�=;�gW��P�l���.<�/���If��ϐ�D�;e����ͷ�f�D��߹�F1��ˋ�=��G��1yl7�`i�Y�w׷������Α�?��~jBF�m���qc4�^��O�y.T�>�SW����h������F�o��Ta�P����oo�}%�~>&��z�7e&d2X+oYZZ��E�zF&l~f?c/F���_=��6���S�<�G��
bBCC3�p+�]C�r���=����@��7$G/��`�8*)�k��ڶu�d�\�!;D�% ,8���g�*� �g:g�'a�NhY�X�l\S���)�,=�P�[G�P�6�PSq��F�����"�QJt>�|�ZLO�A�}�p<`Okl��Μ1ϖo^�N��y6�S��ꭷ{R ��k��S��k��g��kE�M����s�Dmu������Qki�K���N��3nڏj*;S�	��q��ʺ�&O�e�}FhI��5�:�)vSY>Ǻ6=:�}c"-,�Y;(c��gi_H#�qP�[�/���J|4Wx�%��F����NQ�-9�L��-gާ���^ յ2�@iU��}%��M�;��8������;�P��D���D��V��o�JT�o�F>��?���^m�p��G<O��Hm	]�!�\Scۑ���|u��<k":�c�i�+�i�PI䃵����ᬂ�釟[w6�>s8��x3R���D�0Y��m�꧘X�OY�*Fe��D�A�0�dU��ɗ]�:$4�b��h��f![�����=�M;��=����/��Թ�˹|xy��Y=L�����$�[���^c!�<�$F~?kn�z���~s!�e>�q�����:s��p�y��'s㩛qSLS{��Rm�p7t��y�߿�9p/�&S�l͜�Tz��<e�>��09u�+K��_����~������T7m���h��-t(SW���}�:/�!�$���i���B�Ģ6s!Z��-�8��˗���9�n!D{�I��-��mڲ���;&��6ފL/''G\��ئ�x��������!��CPe��
�nd�e�����?z#HC�[񳻻&���-4"BS�:������b��2P��mc֚�Q�����(B$�>n�+}}�̣=oK���������k�"e�0��k��?g���$ւ�D�|rK5y4W{��_%�,�������3_B��8����@��@N��SF������Ҿϭ�!oZl�S�J��n�
f����A[@���6�.��\��g�����^z���o�E֧��#޿�C3�-��W�q43�.۶y+�p���{��#|�m��yA��������83C���{�i�5T�����䝣;g�n[��؀c�B��3�1��-�\�T@h����4�Uj�"O=��>�#�T�r�p��M���sn*�eJ���Ȃ@�BZI\>nf�f����4)6..먾�ܳ�q(�v�2Ҧ?v�T�w����}KT�
������n2�mn~�?���lz=��mEEŒ��,�>��p<�������!�	'�L�Yo0*yINV��64x.�G�f���X�+d7f)u}j7\��\Ӵ u��g�]*N��8�1z�o�k3R
�%����4�=��_��j��<�����yV�����~�[3�ڂBQ�}X�G��	:��fQ�Cb�Hn�C��P��UO��WQ�m:`�4Y���G�.Mr��������Q��O	�V�����e�㮵�*�V��@�F�)�0��縩��A?����Yn�)!�l`���/��c���buԡŵ����_�GƦ����օ6��n&�9���\58��w��Yo��&b`+���������4	Z6Z�����+���� �w(���Wj��\�u��N�������C����{������sԹj/[��:��@��C��t��#��*���pm��1�-�C\��0���쑉�?KF�L4Q�0����>�������4% "re"���d�?����MC�D�A���H�v�#?߃&��{��o;���)�?�fq/���>{���)?a�P�*����Ä13T�^q5@�Og���H1 �zt
���9��MD�A�'C�x�%�mҺ1��ϟ?@��1%�h]�zUbO��g] �A۽"	<{eL�Fs0;������AA>�O@��652�W =�����ɐ�6�o�E8Q����!�mlj�;v�D��M����=��h�<�s7|���͔�����J��=Z�nV��/�h���AO�fgէ���=�����_|��8*���v�xf��`[J�3J��������������������Q)mo�n2$y����qS^%}���@�_[uX�'^>#�j׶]XGٛZy�t�VbkW�]�;EC�Tr��ٹ�� ��P�&��d@;y�OG��f�	����bZ�.	
:�&~lSS~QN�Hek�t����^�
�DV˄� wo�����N���xy�l�lFU}�!t��Yq		���:�,��7 Q�u[�Zr����{����Wr��@vO�m�NF�g�2�5�<� �74��s;w<�@�gn��݃):�GRB���P�9�4��$ pݪ�Ot���M�Q�����Dw���x�K*[�K�O@��S���HG{�m!�K��Ši�?e�xP;O��O�\\��z^�(:L:3ohkk+t�p�b�1,4��Kνw��3������'�?{FFz�����3*�ުyDS{{{��q�<�H~Jc�W���wYXY�/��Q�0�1�z��
fڃ�qD����+����u�*|�jب)MQx�?΂�X���o~$��C�}ra�"Y�it��ׇIDޓ��ah̏�~��ݻ���Û�)L�,��Ϧ�{�l���'x� Y��G�PG�V�CCNJ4`����L~���6��K�T�C:������T���q���	�m�O\�qM|(�yћ��@��̐�N��j�����Ӵ����5�1��f���a���������W��Τ�¯J����a�dW�Ж�Wsp��N� �����+����j���#�L�-,,��P LXOo��o�E>$@�@s]����'�Ḟ�7�����Lt�<K���~��z�ݽt�����r��x��ϺEm����ً��XHZ��ɐj(u�>>F�|�)TV�4&ߟ?~� z����0p�'��۠�����x�f����O�Ő*�t*L����E��k_SP��>���VG^OO�:�����6��v��B�\ �2O�^N�6��*ܮ�gH�682�a�Yd߾}�0�	��ૌғ�M�ǂ����_�45{6.Q^���˷J
+�~���'&N4��ƺ�v�f$���eGGG�C��ʖ����������ѺY8r�����솆�
�k$�l=І��[�B�G����b�q���ܖ�S�N�x��,��~hu||<�_\��:n�ʅ���~M�u/��<�r�R�������乍^�'l.T ���㾺����Rj�Sk� ��t]>6xN穙����պ��<����E��$����	����7B-���ihO;���.�j�	j,'��� �'�hN|��'X�ߌ��������u2�79�k{�p�44�����T�PV; �HB�C��@ͼ))	��!����8�n� %0�8�>7���mj��1wU-�'x�E�X�
3�g!>>���$��L���]p�"/.Ϲj3��ѩ����`�s���bl���5h�K0� ��2�D�L�ی�z����s���)9�%��ڃ��$˵p/Q�,�p��vG�H~`+����>}r@'�t��E����
K�f�M��8�&��8�Q`ٯm�NHB৥�o|-!R� �*�Ȩ�vtT%�rd�ύ}����|��X�����C�̓�P��u����g܄�Ms� ��G^�I?PSS#��	=}y팖�V�F�$&u���G��SS0�@`��lįcO���֨ݺu+ r�l�z���{@�)����:z�����6��eeeZP%Rs[��FйKr�pz�����5�$Ry��QbRSyڛ�gwA����\�S�L����o:��3Pv?���P-w����hhh��d��3۵�����[W�0�V���c��QOlA�8�K��g��FILФ���M(�'��E��*�rrr�����]#c��W�5j,�K|3`�B��ε��>J����̮��k(ml��+�
�����s�p���[��V"��ΡW�
l�b���q���v��,L-C_N,|,u�=�`�\�|<<������z��{7��UUU�:�f.]�́�V����.��R|'tx��dv� 5e>����+=�72�W��S�jfk�������i��x"�.���r��TCC��9�bRf��~��Ĵ���$���>���\��\XX�y����63;[�% �ONzz:w�jFyx�O��G��������h[p�x'��$����Ycff�j�Ę}����q�um��_���N��{vv�G�ٹ(�^��-���c�����~�|������;���ⓓ{����`TB  ��.N��n��yu�;���H�v��qt��=��*��
:����f��C"�2 �h�Li�(7���WTQYd�'7R���BCB��R�v�׌�����F�����07�g��u�0;Q ��5��V2��	t�lm�-��Bb��Ĥ��ʓ�mR��D�X�3�X6��t�u*~*9��.i$��M��,?RUU� �9Hy��+�稨�hN��@/�$��Q��\�,M��#!���yʀ��&L�~�3��?L���{����S<�bU���ʣb`s;�6����W��B�;]P�xKQ�)	���c�kv����m8�}������A�9�V��e� 5�%Tk�8���?ߑ���F{�V�q4s�z]j��!�!T��_.�����a�0�bg�ڷ�2bQĴ�������7y�sҮ����VŏY&ȱ
�U��T��pX������T�]K@ۘa�.`���`L�)�g���'1�����^s.VsO�f�_C��g343k�S91���5_C�m������u�`��Uz�HV�����z�x��+�$��x��w���?�,�#�X���ؖ�JȠtbu�~IHo��F\;s-"�ݻ���Zw30�&�t�O�K��ڼ���(ݹ��?���ջ�@:�a����nkhP�[��	�y�l����=�؛�v���kd%zG$�j����D�9���G���>_��q�
Ŏ��{�HH����;��c�	.��=Y�"�\N�8m�g��WR�A�Ӻ�0S��g@$6���w�X׋�k�#ebb�����痍����>z�}�;m���#��'�YM]�l����Y9�eHcJ����J)+7���Մ���A5f<	B6nx�n��7��ξQ'��v�~���h!нnF5���=��l��B���'�W��i�L�,��Y�ʜ��,��w�
&5]V��Igv�MT�\S�� ���˝챡���S����N1�Ǹ�wEr?�tz��2>�|��By�Wq�]J��MDp�ܪ�����~�����ѥ��dF��U���ӗ> �q���B*��ګ�β�\�;�n��޴�X��L��vG_���?�o�;����v��~���|�\���M.��<���A�����������J��ϿG���4alU�׵��v�O���906�R�&+��Vа�[��6�I2��/��^���^BBV1���n�F���e�AOI��{���:י.:Bp����6��ù���'Ũ���<kg����Ϡ����O
�Az����&{:p���L�7�ZX��rm�3��hC��A���6�7a-y_-Z��\�%&��T��J�֫��~�5�˃�k!`(��$a^}��@��lœ�<]�ݿiΞ�s����-NWgH�?�>�_8.�� �4&�o�� ��������$ r�Z�ʤ�<a�=t�hZl�0���Q4-��M%�(P��EG	�>R�	�m$mggg���f]�t�Q�IO��H�*A�#З�J���:L��P��I�T����bbu��
d�s���٭[0����d�T���Wɮ��1���־/u��a�R�Z;��rd#V-��%��*��Dg=�ͺ�U��'ƕ��D(���R� �),��W��X�&ί��w���
�����Xk"��f�4&,d�A�"r�5��9�H����ݛ<��t 6��.�n�땯���_��'I��H�jq����N�]諨�DGF���M[�����D��Iqt枮e�̲�+%1!A-���kX!ꀸ�{�	¼T����|S��Y*RS]z����M�J���6�:s!fu����ѩ��/��9v�)�]8�t���L���e���7��$��M�FV'��i)T��`���ӅJv�K�V玩�)rt�KA>��a ��r�Z;z�hZ7�Tx2�|�W%��E}#N���2���p;�&EHrZz</��J+5-��u�.:J5걱1�{��w~Z�IWA�"�ozR�W�%�ݻcRRn_�p!S�����ꪪ*taS0��Y�ȣz�/S���̧��QT5�wT��'�E��y���=���mb#%&�7��6�����d����w��s�b�Z49n<��X����(� �łW�'j��
�~��3��mȏ7�cu�Q�, �q�%���q�&r�=�d!Qg�
��&?i٪���F�,%2���#ɚt��D_���[A��PhN��Z�l$�+'�tmҩx�}C��X��@y9��h�(��;P��厪�]T������_�'Ȓ�p���?�~o���$G90;;{�y\�רycYĩ������J�+:OMn�2~��Կ/�� #��F�A��A�ɀ�y ��W9���.$��ʨĖh�!�;���f��K��0T�Y�{�O�[�{��K+��X������gF�o�}���/�Hv�a�.\w}�_G�s�`�:���1%Z�����?�dh@&T���5��H����C�������K���6;C=�*QMu^[�9}������;������x%��'��Wsg�祟>��U=oimM6j���0�t	G#`Ҏ.��z�uC�@��t7�Ws���!�./��t��bl��~8���Z�m2\LL���8\|�qd����{.I��S���tHA��_��ט&������oJ;�P?�0�d���;��B�C���6���N�8��7�b���P����t��NB���B���kM���Ҁ�!���Ǹ�����{q��Qa����e��bH���1	��Gxq�.�=9��} �ސJ���ŉx�V0Pۅo�S
[j���=깾��lC|����/�4�焄���|'�~����@(��@,~�.�����ꄸ�C9&��^ܾ�i|��I����ymW�j7{�n��]��Ŭ;1�y*�����"�]�������|��"3Ur��AV �P/��'����=�m_	C�^��
����3�h�ݐ�=s0N���)ce�$���]Lss�c�𷭭�+�3u:�t��Udee)?�	��-��{ŕ�V�T��Օ yi��<r��5n�wEh@�����a������Y�K�q>��S���@��pLW%�&��Y�H!�,�`�1��1�e+1�z������0W�����ٝ�ͤ�s�ٯ��yK���#.��(xx�`��tp�rU}�]���z��� Ө�Ǿ�N�n����C保Bd�T�v�3r� �^�<�*e�3�3��ֿ�#]�>�O$��@�srK�"��޾8X�г���yE�3Ӱ)8�C���"�GNq~������hw����Gt�C�y��}LLhߔM�E�i�A�.���H�"`� �G�_>n�ϝasY�c��s��ە�0�w���W���Y��;�[��͟����s�*�Wi���Lp���t�4(���i#ło��=
��v|���3 rj�r����"'��g�oW���p0�+Rk]����	u,�
��D諆� d@𲽃X�o��o�c��΂n�Ѻ~���4�+���N�R"�eݎDy��;�9&X��r��C�F����\�'���rRT��}���-=�z��������:�.	�|w�e^#�|�ki�^�_�+��}Ļ}�����:�0�U��n>b��%��~�'��8`�z��q�R�mieu�~k��p��ȩدGԷj�/�VE�Q�����^��z$H����~������\�)�"�Py�]0+^�	�{@)ESö����ǎ�OK=�nD9���Vf��М���X��E����l���u?��Ǣ�ƿ
���|�j�fVTTD7��\(3?$�D�K��SY�LK��H�G�OaѣqC-is]�\���%�{A�݂
񧡩1c\�.ҳ���.ں�A��߫��p�1��F.Kq|����4�^&�<j��&%0��Dı��S��Ggs�����؈/̥���_�v�����;�]�LX܄�>S(SJVgִ�Ǖ���Є�s��m6�x�Z��3ӿ|12��I�gJ�%`hl�T���AnSb�\>�� �F�\�d���K�oP�WݪŊU�Kc0�֖�Բ��zً������v(�Y+&��?��N����L۵�/��0�ݙ�����ycF��O�vz?���hn#�����>==a�m���~AÆ��Jؕ�Q�8����֦�D��R^Q1��D3�ܞ9�ৼ�L���^��g����b(��_w3��4%��MKK;O�i�V��P�s����3KK�.\��2��x�w'�X�*��V%�qb�<=:������~{[��u�+:��)n4ջ��ː�k���B�+������*R�X��\�e[[qa%0�vCKd�/eH1��c�����H	�>cl<Dΰ�
Ω�僱.w��V�;9]� ���,ME°�C�6ﮏ��'QއTU?G埐�/�Ȝ��+\��X��w2����5{����hH`'g\�E���zg��R�ʕ����������+�q����{�`���U��Ѡ���F�k��ms<ވ��a�C�o"�.�l�Aq�����,x������w�ZU��ɣD�b���Kqo�e�Fw�9�A�m.���0�N�e��*tBG��!F�2���c)�0�?�K:Q"��ã��p�8\Z.�XN�h�S�(ݍ���V󠳫��\}����d�5���i�^j0�tk��O�S�ŭ3�a���p����TK��;���|ͱ�P�2�\�̊kpW���U0�Ĳ2n]K�c/p�ى�ۣ����m��z��I���O�ѓ�4eZ{��=��f��"ܱJ��lz��(O����Zև�j]�G��v�mmB\���5>�2X�Uo�D��`5�� '���Ғ������Bw��� ���z����IA��s,������TC��o6R����ʆ+:��<��mY���2I� J���fV8Ǌc�a���}F���;��f���3Hg�]V�mw�[�3첏|��\l�t���w��߿Wo�Ud�������k��?[���Ww��o���G��!��e�ZS*�.�͚��T��	M��u��Hu!k�%F��,!z<fw�Y/��C�0N��imW�b���U��YvLI�~W����ꭣ���?Pi�	A�k(%����;F:D����nQ�;����y��w����r��3s���s���Juuu���  emNXbr�x��ߔY�&j8Z��/lmm��7�����$CI�2�A�|��h��]ώ�kr�Ôp�0�V7��v����c���Q����v�2���`����u{��_E�K��Z���-�}
�7��\>�ÿљ�s�Y4��{� ����!�6ݾ��x�m�2���H@����5�7thAE�c������!�<0�x�4r�2+���/~�|	�W���Cyטx��3���r/���$	�������`���wA�����.b���PX_��n`�!۴S�B��Y���)x��T�]�>���K��⤧����2]���f}��Ye=��Mt[����<-- ����![K!&� ��r���0,���[����W ���.h��M�F��Ѷ���Ty�"X���ҟN��-�*����������a�������sc�-�>�.
�F��[QK@�Ƞ�hŽ��c�Q,r�mu��X�}}]�cî]��8-�8��N��~���i0���L<'y��,��7��RR',����"</��^�S�U��3��uVPT4b�kE+����}��R�۾���O���D����{�AH��~��b
�d4�8�@2�p�!V'::ziQY�x=|�7+�Q�χmP���+�������}��"4cc"d����Z>k��Ge�L���N�n����r����^�z�&��#�\w=�6��a�8O�yĴBES�7U����l�}�"�!��0�W�1�����1�;����P��\��Ґ��򭍗�0�A�U=&���a����Ͱ��/�&��_���ʽy���%��a����
�>U;�d�v�{`��/-P_5uu,e����L>6_������Aae�j��r@e-����~����d5Wn��sc �b���t�b�W�
�c1'�,�ڡEЊm��43\�C�*�[�u�=� hҚ�=���qm/^�W���C��4I�Y��m���n~���<�$ro_�DB@��|I�T[r)w��ۣ������"u�P�X�ӯ�N�g��V�'0���{� ��[\\���l���:��i�E�յ���d�����7��myz��QkK-l�K�*�!����X��6.:�e9����.�G@2z�4�W:��:���ro�c�KY�QQ�u ��0����]�l�?)��r��cȴhUR��#�Ʀ����e�6�\7"�Z>����GZ}a?��o�n��[x�B'ݔ���b�[&/��q&#:J፾��/+��5j����C�?܇LUkO�*W3c?��T!h�P%�7nZ�ry�(\j�(ǣO�)�&��z��{�������s*I���AI�͒&u����Pe�i�m��&�*����<���ɘn�<�$?�
8\|lx�H�n���'2�:~��\�|W����A}��亁�Z�j5[N%�_¤�%���4�����S]dV��� �v����R���KN�W
��R�-qZ�Cݡ�h�8g[�G?ܰ�/���7/�ӑ� P(�M��-7pB�!�u�?>1!G�7�OLL<���os�����}ԁJ:�">?#��x���>᠍y?:9�3�X{!����laz�+P U��7�v�G��l�3��:�Bw��z u�V������I�� )�����T��u1��� ���2}F���4E��Q���Q���~����"ޛX���9H��6� i�<s���%�� ���s���Kh�'Қ�r��J���8|y�ݵ�Q?J��4$��3IѪ����!�6/_C���*sp�O�N�'$$<�e������uH��g�"&(�sP��WW�n����}�	Y4��
�s�0���;e��"���t1�9:��`�0|�֗㇮�Ӈ���;<N�2���m��i{�9�lP�s�Q�3(X��0b�ߵ�]V���P�tE�B~8V���[qFe�5�ѺCb�φ�O
��Z����D����дWgff��Z���;�|�O��شB.�:��=���xm���k9+ʁ3�Ѫ!�T>w�z=�����9�3�lp_�-�A�c[�Pd���79O����W�@W�f���q��0��/=��O�Ѫ[\�۩��GM<�^��F���.Q�G;�b�rY)�����ٌ�㦙I�~�3��U&����=���2��>4�
�}������|�1::j�5�%��c~s�w~~^������ܦ&]������������H��8KFv�pv�i$���MW�M͊��4�O�Rk���x��y(���&������q�����E����֦a|����I��0j�(O<\��^w�t+���l"�7�ݮ=vr�N�22(�{�"_а�?K�񥢴���P�-��0=��ď3߸���Ӈߚ ��~_�;FF���XUh����m\�ɊMA�Y����K��Ǌ�������f��i��4�$�(ʼ/�
��A�W��3����gY����nϾ�mk�'ə�H*0���@������S�?ikc�ڵ"�����Ke�c����� �hr
��߿��P�L��sz���t�{
���Hr�ʈ�T��~�#0&e\��Y��]^��;;���7��~�������_P��/�.:������A�'K-�c�d���AJ�E�Co+�7�y�&!h7�g�1�^Ն',C�u�~��_	��_ܚ��mO���]u�s��sH�����/��s���&�G/�x�՗!��'��R��eNN|O��$6��G�>�����IQ��Y�J	Sӵ����G�`	m��딓�1偭�|��g�h%�Z��)C���X����q�{`��į�.����/cO��գ���!�m�$�۷X�L_ME��HZ�Nn3������M;��(B֟��{u�+,�S�-9��b�~\b1���z����m��� .\�U�<�M�&r��M�w�m�ױ��	��: G ���]�xƘ����l/�揷l�U�]�G�>AXN���Q��Ѐ;9(b�&��-�m�htB��r3B�S�'�A���\�w�v���?0pʪ[�7�a����&TAʨ�(�F�듲F�ҽz�����
�UU!l�N����}���}�kԈ4��7���nk�t����}_7�j�;6;_��*����XX�[Z|q�f�@@�#G�$=S�>a3~��0����L�~�#K�� 	���;��6i��M:7'E�:�n�"HJv�2U�ZV�� -i͞�o��G8_�`�?���? �os)���.��m�W�ڬYka.::��g~�~�U��ǽP�xD��J�����~!������[ɟ|2�7=����ﾼ?9m�C���}�$̼�.fXv���������ս-r�J'����3rl���M��K*ey��X�#)ejR��cS��ί_�q_��7'���$��i�'�3l>Z�1��$Y�ͯ��������G�Ao���|����M_'��K�ʖ��̦����Ș�7���h������Ûc?AZCOO�K��̀ ��%a��6vvz-f�q��F��y1B���"hhF�@^W� �t���#~VH�w������oIU}ܸ�B	&6�퇢���,��Ć*I��.�L9k���Ё�� 
�_L��\�9Z��\�^0��0�3{����B��M�	53���]�v�'����{J_�����
�3$l&�d�γ�^5���;ԩ=yXه1g���.i�����W#��&ߺR�f
��=�#�����S��hS��:(�c�z����k|���p�$F[�\�8��7L��Zg$$��T%�;���!2��(m��a���iA����o�zqk:*�I3RQ�f�I�0�>䳆�zY�Ȱ��Y�C�O��>�]?= �[�3�ܐ�(rl;����~���z�n�A�n+|���`b�� � ��?M2Y�_"�7Ra3��&�dr٥a�]g��h�[znJJJ����7MO��TJm.����h�$������e��@H{��[S��\�\�8���l�̂��wl:]��Uu�__�9CJ\�}����.�9�)�f�ŏ.&&E�Z���]��]��?*�0AK��+\z\���E��a�0n��1�����X�ǖ� )7��rC��������(�fLH�'�-w�M2��
�,Ѩ�.뻬�'چ'�y��Xz±��L/>7��3�&ȷi�5����yʗ�4!����c�!4��z/7�O�V9��K�����߾�%�����2پQYI�ׂ�g+�b�lr��/�#K��v"~��*$���i%�3%�*t:�[���Y�\�݆U���ָJ�BrD�\b=N#��b|�Iz'�"�τl�I}vXfIm Qo�pL
ҡ��@BBC9Z[oC�u?��7/Ê}�~��~��v^�?��&��ς%�;�F����a���/޴-\ʇX�5��a���ӧʚ�߷��u:���ݝ�'���� 8���W�^��Mq�δ�	�NnN.0X�WOYr����d#q0q��'6��|-d.����>�U����8<L�E1�[_wFǔLjv�Js�Kܳ�w�����pn����<��V���7褓��F,������wl�sk��3��9��VT�\�u���smoQ%��W�~�;�v���ٳ}��u���hyغ�S�#��Ȑ,�8����F�[��.�jK][ډ�"��@�7��-f�ah�/%�h���斖������}�/���f�d	].�[�27Gb�8̡��I-���}�$��X���e�H'�2e�NY�m����1t����^IP�th��$[��~E��etzqw��RӿaMڸۜKJG�W��[�u����T"$����<z�V�)z�Ns@(�*�0Fr����f���s<AB��PQ|rr�t��f���+@�>��[�3)ʢ`�S�C�d��fOb������{�}}}���4ٺzo�����7�2��%�޷_�ɹd�����$��h��E��g�o�Q�/���?�X��H���u@)O�<���^m##cs��"ܶ���^�������]�-��w�8f7d$S�%J V+?��)}�vwۺ��V�,�Z�����G�~���>H�DS����زކ8H+�Y�!�r\�j�3� {�3@8�Gh�(m���m(p����Zʬ��ȩ�l�*�J?��Nac-Z/Ts�D<��s�=����0�\�۬Ө��ӯ3*��.��09�z$�\<|��0X�Ar�����\���z��t������*q����j�j8��� �D��s;a��C��S���\�����%����e�5i�5����h��ܱ���<^������E��.%�#m*��wɘ�0���p�-����f4���]m���*�HSj��k�����H��}��ZQa�v��%Q����*�k���=��d�)-��8�|xshI"c]kL�R4�0Q5��i��2�Wn�w��W0%kƦ��܂����sA���;������'�v��[���|�-�X��N#LRSAH�l� ӥ�VX�����7���Mޘ(�J�˪I<�=}:�5R���<��2�\Ğ�zU��V�<;�ڛ��4� C��uZ~�K���:4<��Ca
o� ��[Ty�6{�^�S��}�/��.*UW/�����0���Sew��~�D����/_^@z�)�Q#"#��_B�%:Q��p����_�nw���O�?.��&hr?�f����Ar?qa*0�Ї�|U���=M�"��?�E`N�����>�)�c��I\i_��V��oy���B͙['��_�T�#�G�+xM��g?�<eG*ϣy�5����e?��6���_t�݆���}�z�$�m�'���8���c�~��
}��n��#��q�z��ȅ��;{ꬭЍ/��WK�&�����(f�Pjd��ݣ��jk�l�
`'Ҝ�����J1z�K��x36r�/9k%l�ƅ	{��!5�Q���M!!a�V�Q�щR���V���1���d�E������%���Bf��$͢��K����F��5��������_�h5�,��Z]]嗕�

sp~��1�\���tИ"�n�=�Y{�!P�����&�OZ'���a�}\|� �@B���L��W��.���Ϊq�?1���c7]���LS6��,e��fMU={�L e��ڂ'��)���[p��#�hg9�h��z�0�W��ZWjL���`�����q�@���g+��V��5 �b��� �:�U� =�W�\��Od���Ba�h�ToǂD�IO�n�^�d�����{҉?b;�&O�	�3tz�uXh4����o�*9ss����� ؔ�������d��B3�T�6��-,��ѥ,��P`�+++_y��x����g�܈	[j�:>�I�}���)��������87'/��`ӭ���j Cǭy�z�EJ���2&,�"''>F�E�����}��m��R-���w��ӈA����ܕ
l����l�Fۖ�d�?�|�)C�_A�����?� v��ߢ�9Y
�����R�:���~�n۾Xl����gZ!՛��������e?Il/���i�����=
3�?}7���X�!F��b�ѥZ$4��Rk�OD=$�vи��U�}g��~����j��'���5B����V�b��h!]���򅅅2����R0�:�������F�J�nάp�y�@�7��̉���G���L];��/~�EײEu"Ve9�@C�!#'�3�E	�C�Z)A�d�����8���Mq�d�q�c&ܚ�#���a�����>�0�� |�x��4�o��a�A0`�eD������u�
�܌>.�ԉi~_o�����v�AL,	�'4��F�[���l�
Lj�X6E.�T�@h���� $
��n9��3����(���#Xy��I^(��,��������3�E��d����;6~�K�k��P&�����p�[� �J��m	�/E��NOk�n����
�c0S�i�m=�b(��!������t~ʶ.���eo�)��sj$���R�p���e}O��Q�����M?P%�ՎK����e�4lrx���N{ڀf��)����#�l���fY!���&���T$��X(��Jb���R�(F���yf��x�b?�غzZ'����F=d�=pi,}���@j^C�L})S,� ��5���bhG'<�u��Q��#��п������~R�-]ː�{�:��F��^��'C�B������ͦ�-J���y�,����&�6�D�����?�jc�΃�.�F�B�҂���^g�v��S
:��F���3Ј���"t�55�띌��<e@醆Ry廫�����f
j�Ʀҭ���-�T�{����#��WؠSjDDDeHHH꿡L���뻱�T����5f���-"w!��W�I@�J4`��O��Q=c�%D�k���WV��k�Bb�(����˃��=E�8�K
�f���
�S�q��-I*��l_����ȹ�t�![����q�~�P\_na\�Cqe
ԍ����! :�_?]M�ȭ?� ��n���?	D2w����l��,m���]JP���i]��2lC�
V�V�g���n}jr��]����"oh����Z�j�`�h"b�����f��Y��^a��i���͛7_E<�a��-�:�Կ���҅�x�u߶���-�������i۹DsWT���{Ci*���~3��U>x��" �2A�������V���7�R�.H��O�P�@�akx�F������ϼ/6¢��(�0�9�>�hx�?��ۃ��1絜t�����g>��_�ꗿ�?��!����@��i4���d|���lu��rRd�Y�uG�u�M�8À�ak���^Ӕ���_����]��M�;��p�A#PXj��xxZa#I���<�.������Ic��w��rr�i�G�v#|9�̜v*ފm5��L�*�׏�{f/�J !|����|�	��-�����>u��緉�22&���*E��%X^-����'�=�Ė�4��e����}�IIIi{����k�f>56BF����m����Af��kl����U��O���4����?�y���cIe%�\�ch��s`b���X�>����;�u�t<S��yg�TX�*e�-����1�(�Q�z�k5��l~ҲEQ�j}�,��GR��S���Rv���J�W{����J������Q�S}�S��쀈*��-[�x.%�Q �v ��;���/%s�����8�@[���:�M����"�Y��6�Mp�"^IG�V����k�n�'���t.�����%F���42P��KH<�M���`�$H�
l�����>��ҳ�H�qf�+#��Ֆ����@�:�����"���Pa> ��)�h44�\b��^qp�ZYկ��/HflV�R������`�#l���1@Q�ۜ���7c����L���9�&a��\���^�w���g��L{iQ�K��A]�E#��3ϼy��U�y�v���<=��:s�Qr�(
�6Zä�.�O�Z >V5̊������ ��}f��N�♏�"���k�)'���\��lH�R�!-ok��@t�����D�ݢ���D����eC�j,�<h
�)L���5\y)�Ho���b�\/	���Þ�e`c�
D�!J_qc��洣3�oA"c���@UZZڗ�����rI��Q��Ԛ�K���dx<CG��Ɵ����������}�b�� ����OKG�v^�7�ncgםĦ;<�GN�2���W@�z[�y�|:+[MZ���36�h��~�E�=rWE��c׶0�dS�NI7���qkrb�)~�BS���w���ޤ���0ӎi>�B��Q���0��1�;ie���2��S��Ӽ@�A�,F�Hz�ΠU���$5���gЌ�($&u�����^x���0�kNi�8�4%�05���s�/��1�����%��ߘ�9RzȖ��r��wf�dN`���A�$ � $����c����w�L�l����_�c��ǟ���ή�@麰/����z#���-:::�rYjF4�%c#f׻�dg?�B����&��J��)p ۰�:;T#�o�v5I�Z��hO܀���������'T���c[&������Is{����g���4�ǘ�7[]��EP����uj�|�E��K�}���U�3_����͠y$�Y(J&8<G�smpQ$8~��">Q�v�D�t(�g��11b�����'��G��� 1x]\�}����A�N�Y�fx8�`�Q
��������UG��tk�sh��P���L���I>zq������H�9�8#��: �b n�=��*u��ߣ��Y_2|���H�p�v ��WG� �Q �����_�i���B4�$��mfwoo[_V�#��Wu�B2�!=���S��Q��j��a�#���9\G�wYfH�����]������/�+��%��Z6Q'���S*l���I���h�V�[(�˻W��[H�H�_�ی��QkSyy9y(���"�]�Ӄ֯��ՑϞ�K�}W�&u/qQtvsg�분)�r ���F
�/@��9�P�&��L�Ǟ��`�[�s8@.۵�� y�tdJ��<e͊W4���:��-@���l����r��lM��q��]�ީ����� ~�.��b?c�յ���rJh:$	��'��y:�&"B���,"L�M�0��=��=�gl#^�(uv��XSQ�����X�s|��S[�	wo4���c��X/�*؇2Zbw��9�f�2B5���[�/E�}�8e���+���������}������E:���f���4��.��/Q[�4֭�����C�9E�����K�ab�2H#=H-⇨B�h ��	6�g��1V�V�['\@*4L]ӑ���r�7�j�\ՀT�NGj�O��&@���k����i�'?�Z���B�{��=e�|��YV�[�	П�`SF�GBqoò��i�jk/��*�����@��礤��zzzԉ�/!����j"�uo��#kO�����
������911�X\R���;{Dvи[�����2''��xa��.��EW������7�hx3%�����!x@(�r�j@���j��J��ZT]FG�Fi�t���/w�b�i~��O*�����Jw�=�hG{����Y�Ͻ�u/��u_	���"�L��ފ��oz���J����O�����:�<��{x����7�Sō�-���&
�Z�>���3d!.�\�&�5̯`���o�lS�6�E��0�PI�v/Id�D��4�cϗEId����u��sf�m�*&J�Z$�oP��k�|{NFv���'������ zn!���"vc��GK��,�s.`Lp�V��g��Mp'�hxy�ⷶ�� �яFH@�L��
3��H�=�� 7���e��dL��o-H���K�DIT�=k$h�h�L�������I�ys1J i�{��f�������8�������L�`d`iMxԗ�+-�����1���	�`ʴ8���.�T� -꯰r��Y�ܻ,4QN�_���=p"l�������z��8�E8�Z�,
�r~i���I�'�����;���ˁO��*;j�eї�^Z8���	���}�-�L�<�D����a#�f`oE�;�������GDȫ%p"���f�؛A�c��X���3����� Ӆ����	�AJ���h������"��ww߾|��9b<k���ߛ�� $\��2�5��I�T�&4�)��׸��/�ß��1�d�ќ���?3�n�fN��gU�<����_}A�*��y�3�<�	k۸�׋�첈���{�v�b��џ�Fw�"�EY[l20��t��.�Ms���N3���$���Գ���Y�/1U�1 }1�gl=	�汩�s_�EjKEF��H_�p].�k��_��/��VC��#9�G����?wbH���.G&���"[MD^_?=��p�+((hj�Ϸ.��Pr�P>��sP��@4\#�X�+(�fd`�v�@z��qfgfFh��w�&H��v����]���?sc���`���������NYi���*�J-Vx-���H�k�NF�]��E㈊�*L>u'/|ӟ����'�4Y�z��n�4ޚ$���I�����3偀�}Gʰ}.*  P��� �����+���p���|H<%Q���d��Ha5��"�s�C�F�fX�	��-ݓ�^�#*��=���m�jA{B���a���������MC�_mD��F�Ksma4$�k�Rnd���A�Ń%p�d���F�Gw�����q�Eq�?�_�Eu����hZ/F��W{��-*e׋=m33��q͛:Iz �츸�@[t)�"d�&)ݚ�=O���-�X�8���<���Z�F�MIM�0�����B��:k�l��'{��82�,�%��Ñ��Ri7���Ņ��+$��גr��ψ�/�'2>�/����VDQ�^���*b���
r�q|�6��![m� t�dhr�:��h���XKǏ ���B*��f� Δ:;<�͝�N�`
9�,�O�� ���N�?`��2zC��㊬Y�~�QȻ廙;}�?�$� .z�@,	��-��u䝆��$�w����"�i#9�Ej��888�J����8�-՟>=137w�g���
q?���1N�ߧv#www��Y�.[�V1��Bᇩ�$�o�������Y�����8]kO����P�[ʇ�Y�C\Pk�w��+�p�<�M��)��X�B�hv2M�l-m�7
�m���nnM4�9���X����^vC�v��o�VG��-�2=�:��	���K�_Ҿ$>�@*­��ÉY��ds�J{z�����5Е��v
(�f1r���?�<t;n���2Z�	���a��c�S��H��9*�8��_�v'�@���o1h+jh��� �ypL�PB���~�J~w���-2���D�s�k���>}j|wu��_�|QŌ���B��zY*w�=��S���Ժ�41x��� ��\��S򯮫��,
[2r_G؛�"P�#�m=�|�=�r �p��9Ą0�� ?:��5�'������m��cf���|�Ȟ٧���bGF��{K�
t'\���M$���23��2��H����2-4��(�9|�����|�F	`1���M���˼��~Wj[�W��k(A�f��f?[-!�a�bc�F�壸��?M��&�wO�+��\\.N�9��xT��_i�-���[��B����'8*LNZ�(� fӡı���OΞ !����
q������n�22��B��;�c��|��#��m��L�� �jj29��jjc�Ilk�3SF�F�����.QNd�\$����6<?`*l>�O&N�|͔`�+K����YH��p_�ݜ��ZddW1�M���$��~�猅��)[��y�����M�\�@1��� �: �9�O�wǓ�dCqM�A�h<nV�x� �x~����y��~e$�_�Ǔ�������ϼA��~�����]kl]�+ W9+��=���+���者��9�Q��i�,��h�w��ʾ<�����E¹&iu�������*ƛ�]ԧ�lV�rq*��KZ��ו��$��]�w�����y@ˆ]E�b��9mӬol��찺�
����A��n|jj�����F1�������)|�2��K;+��(��̄�5���O���%EhA�����s��l����;Y�+����lM��Ͷ�n�>fJ����|>ˁ|I2e����ݙ����3��?K��|߽����>[�O.o�k׎"�W�B��F'���0<9�*��)}����3�x�����-��i�'f�&1�sχFM[��������:��A���n��qx�)}�K�{�6���,�KE>����bps�kG�I���weҾy�?���($D���*�Xb����Y�?��Юc� �>�
�0D��GtJ.V���o��輷`��-�gA
�,�\7��ۀ2p�Q-���r�gd�����X�	��	RDs�j9����VY�%�9be����U<�}e}IrE���d��Ɛ�>�h*����:�/vB�z�����#�N�o���[Pr���OѳI��8RS�g����~{����A���G��G*/q��ُ�%�V ��=>�$w��8���_���\2�cO��G�:�q�Z��;�r�8�C+�����T^@��	�s�l�]I,����-R����_}���ܛ0�=9J��[��y��w)�N�f��L���3�M�=��F�r��d���8}����o+��Կ�i�M�Hb��M�c{���c .p������YYY��q~(�UZ�+��u��09<�*����϶�daS���CBB��������C�)�����.�����e���dQ^�_�����"  �g��m\D+��_�=���f��X���a��=��
/�,$����5��5��^�����^���ش�z�"����C	���2�Zj���7%�S�њ5x�BQ�vW,~Z쐍F)Y�՘���t��S!��d�{����]���e\Y�����D�B_n�����۠���+�]���U7�l�?U��%�{G12a7�������R�V��ϑ`���L�f�:�u1��&��o�94n3 ��FB�ѱC�P;�x�NSRRj�)��᧓fm���\gĳ�C��;�;99��{�J�ݞ��ߤ7���3[m�t�ď�?M��ШI8�V���uYY98�s����w�e��<��h��[�$�T�⭳��]yxxEz�/�ӧO�63s)c�R22(�-<T�{��^�Ō-#�ft-[�T�*L��ӂ��>環%�0�=�!�~]�~g�c�f���i�ܣbo��Hؕ���aiۛ��K�F~ k����G4ʲY-K�Rgvz�6�8��yN��	�+)us�͝�ö[�Ei�A_��>�Дh�q�1��r��[�S?wƩ(�.t�� �����]�^�8�'e���Č"j�I�uWLrD|�PÏ�D���$ �&8��B���৯~����oVI�K�j&ͱB��Ds7)�R� ~̸��ߟ"B¨��S�	�mXcB{{���$ߙ����<Z�t�1|�A���#��|,c�X�@9����od׆�H!x�r�.o���8W�[��J�	�> ��Ru�P+ޔE��R����u���m�`��h"B��-��R��� �%%k�D���&�Q�!j�3�����v�T���Pճ��l�$Ѽ�ZHL�h������.郾:�r.?��.�G��tw6��t"2_�B	��ow���ۜ�W~=�,�h��+���M�H������ĥ����`я�����p���i"���o�mo=���-�-�p�_�D�5j6�D5��f�})�,�} �Z��ߪԃ8�ی���2z�Ɵ����,Z@Ԫ���ҡ��Cn�tTb����8�G�H4~~~�@��.ќ�����8ۭ��Q�ۂhDdd�㒘 Es�aЎY���in��H��' ����4�P'0�!��Ws9��U�^q"A�����a�Â���"�B�U)Pg&@��D�W/|�(OX�Z@�ά�U&M�@Q�dR9o���K�8$eo��� �}��YK'���aP��U}�b�'y����L6������;!�v1�ݠC��t�^�R^����չ�JQi�g�:��=�'}�п��Pn�nB⧷����'���P����M��ʝ��Fy"g�De�9t��>�,� �I?��_��-���c�h�{�����-ܡ9A�kA�����l�E�U���Av�v(����� kp�/3?�A�`iaOѓ�����"�ǄK�d�"��&H���3��eϯ�+�U.�>�"�B�ܵ�t�J�.W�����C�b�WO���I�'�%��E;*Q2�?4�>�D눋�>�F���ES�G���H��*Ƀ�F���4�~&�(�.���;]�Hmǟ
�����,@�Ӹ>�Y�৻(9�.==�s��7�-%꽮%"�p"��ny��쏉��%��o�=�X�@�d�� �t�7ՠ�&�E�Tid���x��N�;dS�|;D)��8��9nf_%�'���7<�!:�/ �fp���2�0_�B/$�W�Y���مσz<�FK�'�B5�`�1�~�"Q �)�$a�8��Z��g��':%�0�X��;���+(H�`��F}�X����롗�����!z.<����Fp�,��w����jk��joA��za$6�^O��g�^�����G����ԦHhC�t�Q�'Y#���(.Zچ
>�/5Gﴣ��m�O��-6�q��W�E%�S�!�.s��Z(���N��?m��B�w��ڋ��%�j���/y%y��BTgH��ڶv���K�_�r�I����l5%�l��U��s���Jn��z�������6������{���#�ÿ�A>=C(,,TQSQʇ?��2�5�0�<Xt��^*�y�6�'�jE{��H������Y���\��T<�-�,c��zG�p����<�,D�x���ӎ��gu�R.���ٺ�$a����+��,�[�>H�,��<ӹ�`+�o�8�`(�	=Z�������4w�X��Z���B�ʨ��9u*���R�τ��4��<��5]KQ\������<�rQ����)؛������?�רp3.�Ӿk��=j6��t��j]U財��;�%l�u�t�w)�M�i��RS4/���$ɟ���X̶�Ø�J�$��O_�/�dA������T^�	���|�+\�����c9Bv?y�9��,�;�}�2-z���YxZ666 څ��~���r~m�ߒ��@��1�,S�#"�Y67~d�Ж���'�ߧ�:���0�L�d\�����iӖ�Z�ӹvtq����2�E������-��Ԥ�h�|Z �a'�3����Y�#+����*ֆg���B�G���*ݼ�,_Ms���u���n�5w�w}�tm|�����_D�kz�4\4=����JZ���`�_���C��$����$�P싃���K�����ފ�W��R�_#��z��nymln҉�REJ�Y[0cj_А���)���d0( 9������n%:H�o�~���3�>��x�륟���F3-��Ĵh�t�����/DXhI�29���l׾�cd &<�̱�3����P��W�Yﷰ�Ÿ��j�myu�Yr��Z\.��ĺ�Z~Uf%��D�T�����]o�����T�#}�����vH�|	���:u=��H��&�q��*���M�1�'tst���['�"<����я����x�]����qo���m4��`~��Zy����L�;�>����%�`�IPj�9n,N�ml��D:<�c��,��ڨ�>6�լ����y� *g� �,NQ�/���*Q���@m��R�N�M�8;J���m>��0}�W�3���!2nn������XT�F����sE���v0b�p�R�>���Κ�x(}�X���7�w��2��u��;��A鲰z;,F��F����j> n����%���o���}��N^��F��P�5��<]~{VG���kjF@i�1�ٍ?�bK��2���/*���A���$��@��	��Ѥ2J�?��#+޻����B�#s����JF{�<[�����]Z�p��qR�p�Y�p�3�dL'�G���^�m���7G��T2d*D8�"�~H���X��Mlֳ����_O��|�]s�ͨ]��V4������	�+�*Yn�!�q��`s�ѯ���h��ӭާTR��s*��>K	�k����p{y��?]��؟����|�a�/�@�uvJh�hv����p��J�ptZ��537?Fbǭ�q�bR�A����y�oT�ޙ &1�}�`?��M��W'��G:�ͬ��Ȉ6;��p#,"H��:{��O����Q-���<��!����8�8��^�ϻ��\��1�����<���V24V�bW�=^@���/9u���_	
�15:D^�,I�q�V0����ꨨ���AQ)I	�����T���DABZ�[@D$��n��x������t�q������8����,���VՓ�%>?#j���f�wW���gz�?���ܒ�Q�%)S����I4p���g���Y�8)���z��M�5�*��[1����t��ӕ<�qG����ɡ��Ɔ�����<ڛ7w#�Eԕ��A���B�8����N(�*��z����~��R�Yn6H����:��Ɗ�b�'�	fo@`���3�C�X�'ƀ�d�r�c��09{
���m�Ņ���g�L"5���4��F��\J������LcH�RD��<Jz��Y���+���a�Q�>Ɍ�s�v .��]F2�䔥���=�9�MLđn��[�W�Y��u�/IZ��7����ܝ)�$���g����V�q�C�w^�Ȕ����`ëB����&��)n�3A[�;a%qڈRΆ�����_R�3��ӏii}dc"�Ԓ����ev�bC��@�)(Ȗ���$���P<����M���0k�j_K(w���2�8�G O;�O��Ut8��U�|-b(���������]_��~s�����dm� �u�3�);���`�n��~����`����##GMMa����&�fP6ٴ�z���4>�C�6��o�q��Ȼ񒯗q,�@��Ri�q��"�s'�����l0d!��!沅��*;�T�ę�t�t��Zf��[p�3���P������b�xxw�%��7������e��@g�|=c府�@?�N�������}��*;�v*-5��Y�o�.�#Ra)���q�����у~mzb��|�8T�{����#��:)	��6{i�ƀ7� �#���(Bʱ[Uuik�3%ẍ́���c�)�q?��p�0�c-�a���!�3����g��k�P8C�B���eC��-���RE�58�����q��ʓ��c���'��(
>�̝A\"���@.��^�4bm͔6��nԎ-<��n�&�䟺��A�"�G/���.ICq=)ᙢЧT�M\;}E��x��+ؠ&L�|}u>�n���#���v<V*D�N	6_��?�i	K���"�1����5���J���'K~T]!�׾���[}�ر~yz>���8 ��8a��V+M���;Wơ�`�U*)�ZJ@v9�K���E/��(F����q��߷"[��/k�̲U<��k|`��س58ʕ���+o��>��\�@G�$��f�;^ցR���_r�}W�*�Q�K%��v�Fww�}<<?_X�h����.���T�I��3s�(Kt|dm��a=u�Q���x������L|����"�k3�&b���U�F󡷣l��î�2������",���3��ln^����K�/�Φ�,C
�`?8kwՉ����~�g�̽�Q"�^��%<&�d��u3-�L�h*���<��U��o�@���i�r�%���:� �^�����4���9�f5!�L�|Q��l�-�O�Zr�y]{+s�ߠ5��"Lj��a=I��<<O��/��T�� ���D"�65��JK;��?&$�I��y�R1n��������J쩣z�G����m1��r�I$0L����Y���̺�=���+��d$�A |у���-��*""�l?��`[��X0d��j?(iw^[yn'P����)u�_v��UX��u�����6O	�5�]�����������	��Esu����^q�2�'3O��+A~�*lGԳh�9%���4�?��R�$����FJ�#�a�>ߔ�U��L
��#/*�~�pn�3I|,,�2�--�G��9_�ES���ݷ)j��Ds���gTÍ�[��v��x��:���T�@�k6R�Xϣ�Q��%&����]�hʲ7�(�!N!���N�z��=�������x:!����v�Q��C֝m�<���|Th��l�wkw����;����n��G SA�]��}^�.Ш����-L�����A�0��!�ى��S�z�oEruT��;g��װ)�?��)f9Y}��e�C�)A��qbbb�ϵ7�*�N�Q�����������$�ת��k�H%]�F�j��&/Skk�7����X��PX��l�0(Ƹ��^���^�W��p�i)�ܢǖ˭;�2�&�vߘ2�K���9~�8h���JF؍�>N`gWV��['���6M p.ۨ�
�ZT�$l���q�멉dm�[�!5��s�vME��M���b��ɡ[�Tp������X�Wҹ,���,�i�;3���T�C����e�G�=���8~���HL�hA~~�H�6���_��Se���v;0^;r1SD�o�����f���K�n������NX��!,��UN��O�^{k��>�uT'��c��y��r�^d��w��;f/"�B�f�l)*�g��΂��[~�z��[_��Q�,F]��PԷ������5'=��e�N�M���y7�j�����p$zq��R�,�߲�iXG���	� ���/�ҡ�"�H��?(����Mt��*��/_:��߯U����A.�����Ee�g_a777	yyq'��5b���(���J��?V^r�u&���[7��m��o���Ӡ���`�{���~;�w��
S�r��ul�S�s����7+�÷�a�xt�t�n�(5��f�vx��.�{; ���*ϣ=G�}�~�#���&1-o�����o����9��x7���鷯e�p�_LceKQ��lw(�x/�Y�oߖ���`��1����5�z8�-6�Mߋ�$
��Xd�P��9u��hck8e-��n���ь��K#�w���G�ʧo�'h��{��%%�t�����Q`���*E���F�
f�Hrr@U�G�;��� _�b��֖�@+b�����p�>8Vi�+%%5���r�%��ʦmV��5e-�a�#a�p�lX/	%�ZT�������ie8m���ۼ5l��ƅ�d�[������o��	�ʘ��-���BTz�0���M_��f����if"]���h$p���oK]7y��*^D��ś�xE�E��x0���:����5��O�:"6>��6����߉,!	�n�D���`?6v�6�m,P�����Q^�'KS�����ЇJ���l���������[X��b�~�Z��E�D���y�����B]��m��9��/X�B��[���l����H���̢�
V�n{��R�R��̒j�1aI*1�<�d���ckw� �I�j�c"^�/�k����_JJ�ux���~�҈If��O���J�A� &�O9�<J2&�`�i�ܸ���-ѣ��U}r�w����Ty��<m��y-���]�gP&@6�>P'��劎�x2�^���C2���/��6M�ڏ��"��Ԁ�:f�%��p'�Z�@�Q�>#�u��#�Q����~!�i_��i�:C��E��51t3�2�o�/j�f�lx'�e�N�Y˒�}����i{���CSS�	K�|(O�3�w��*�
y�N��OM��k�~���z��a�ٓdJ+@_�0�ى =T�Z����tGd���ng#�LrVgA�����Wl��B�T�]�^;;s@]�=Q~�X~r��rX��I�zM��-��� (�uԄn�z�a����ù�MW�p��e'
w���ҽ)}LG'@���.�
 �2��\�=;h���)�U���?�z��"����i-)n<�=V5�%�a���ܐ?�'q{U>bVvh�H{�k���"�;�����W3���B"��t~��G���slg��{P��N�#  ���i�KLr#��䠤����S�۞�����P"�KbNNN`�+=I܎4���Ӿx���2�U9(��QPP�Q����`��R�5��i��\(yU��a����ߋ�w�6�����B���\������}~.��e�p�-�58x"&[1R�W��RPI���Ly�v�!2�nj�}�l�5F�07=J#T�\.Uכ��R��*���%=$���sM���iO8s>�Ѵ��������S#���F�6w���{��q�6(��@�X���k4MMM�*��ܖ����L

��"�����&�~>�
�1n�W�-s?2&%�͙�":b��_�r�L?�I}�b�>���~Q�3�v``���F�E��t&Y8��1^��	��D�!���g+2×�U�n]]M��j�A%X<�v��^{xEw��&>��5=��1��BLd��Y�O�[��@I��ӈ �C���fI��?~�n3��_5`��M����d�^#���vF$����!'V�[���쌸Zz���X&&qKw,CTJJ�e��T�===\j�Z�8-�B�DD����p5"����;	_�@�z�0z�~�`�A��)[X��?��$����^�bD��QѦ��X�\��J�TQ2[e��F滗�G�ܳ}Z����g�i6r{c;���\UG^�L�0:��IT��l��o� ���}�2������>S+�.ʲwE�$�!\@0o0����6/�v���)�'�c6�O�z��17��餅��L�ފm�%d����CEš�{��h�*��f����1]v"g��K��j�$r���/��e��"
z]6��&i��JCi}A�T�Z� �u�D�ah�}���|G1������%�vK�iߠr����cF��00r�8���M�Y�?_'*#�2_K�jG���S��&��q��[�DC�m6�U1��/�����JYo��w<���3� ��������J����u�v�C6�.�(k�6f�"����|�C�!g���ǰ��O8��W���3�qc$a�Q�<q�����0�N#�o�㙮��|6Q�}�k�b���f��Q�ר%ϻ�:�>�j(4`�[Xx=+>u�WH��d-Ȗ����K��������o��6P�?��PUR��:Hs?_�U��*�����=}p���u?$��e5�^C��~ ]�^D3�nDCt�ӱ�H�@���zY�J�o��0�����}���I�!�Ϭ�q�Zܦ
T�)���&5;֤�+������z�Nr����G擔�
�(=$l����7���VWQ!����ٲ)8��M����a\5�AUfV�co&�.-P��lQ�h�������X��w�,���������*�E���j-��7�V
iZZ����rY����6���ݻ��xߙϡF��E\x�Ul��D�`*�I���SrV���YVb��T�G=d���%��:��xÖ�F$�0���1mZ�u�v�8S�	�-[��c���ԝ�\��SЍ���U���J�X��|�DG��bS�k�u����P�\dǬ޳t}@Vg=f�7�Q�7�Ф���q�T���tzAȵ��g�Jh.�)Q��y?�"*ؓ?����n)�L��%%{���3�뵟?����Xm3˔��Q��C�1�f��N��o'�iboik�%����'�an>9s����n稈\��w<Y"���F��	!��l.��Wg�C(�򜒅ٶuK�:Jbh'�X�3�ޅ�$�+?Ϳ+64�͜8�G+U����x���i������Y7��EP*s9եz��M���l쪚n�\�o%��=�@Oy���Ҧ��EC'C�����RQ��xLRL�e�ӋL�!s0yD��*�\�\���-Ӷr�`�����u�aH���,ӧ��^U[��GUU#�lB��=|M6"U/��j��'�H~E���t�����[Io����� ��3e+(*zѽ}�����j���OUuu{Љ_g��{ނ'~�sIS��J�L������DfXEQ&v�-mA7Q�Y7�@Lگ���}��ݟ��'�e*�m"�� ��o�̊
���^G����_����7�����_T#и���k���kQ(��i��w�z:��$����]���hq�j�j~�C�(^N�!�7Í��vx�q`!��/��T��[%�_?T�����rP��r��q�E�l)`�ƍ�5)),���ЗA�)�o֫w�RRV��!w�r�NX�C9VP[AA���jltt4��oB�T^��2;�Ah��?����}��I�N�]#(KS�����X�/C�z�źd�e��P)��#�]��{V�_�`nƣ��u↤�ݙ�����u9���N^�wihZ}�����NӹreP��k�A�BE2�{e9��DkfB�7=�/�Ӿ
j(e�|/���l�v���2ő��KT8q���gS]kX�>3�����g�X9L#�/+��C_�\e�5��!��EH9WNUH�ω[AZ:���[�nu5���'�7t�%�_�]]]D�Բ�Y�J�.y������ T���XAg�����ݜW�U�i�coG�H67!_��v»?J�Q���hM�e~I������{�˂"��>�~�=g�H��j��Fas����1`a��,N�
T�7�P!	}3��]���b&1�Y���sם���]�Ɏ����8�����JCNIzr��ȕ��j_9Wf����������x��8#�C��tԮ�d��ǰo��Ǚ���2��$4�����
k�j�Ԣ���Y8%QD��I!<###s�e{.�[.��ӡ/gUQS����}y�A&дӺeo7����:1�5<2�����I���O�Jw
��3�[�Z�,M�)��=6ֶ]V!C���+��?��Ӟ[J�n�G>�gS�=6e�^w�=��͑��Gi!C�6�s�G��W4�6�J3��*�tF���d-F&}�����;%�U�J}�3XTiS��a@8y5V3<�cH�H��Uy����ƽz��j]#-���6�u2�FƂB���ק�j��چ9��d��jj�X���ӟ)~r����T�xO����˫��S���^`��M����h��r9g=?a����b����e���cP[㽮��~��$|���1��Hv�%LO?��}��A0T�Y��ьs�5�*y#�'�,����$�`��#�(}���gSV�z�ޙ��Y�n�H����on��7b�Tj��}��S���dy�t��9�g��`?m
�+�+�@u�S20��˩�Iސ�jaYޣZ�|�})ǃd}�B^gD����j��}4 č���1
�/Jq�;���o�^,��ri�'�
 b7�	�I���{�Y\,�W�~��=sSS0�wqM`0�-�+=vu��]0d<�<-Z>�wQ��.9�����y�=^��vC�0�zp�/�F�iφ>�V&s5���`m��V#��Qj��A����3��M�g��M8��_�Ṡ�9�PO���~��-�Ƹp1ʉ��ҍ$٧ �z�ۼA����7 ]]֨�i�?����SW���r=�Gn����<�d\�ڊ�1=;��c��r"������=V.lffFOO����u����yͤ	�u@�v�����R�Ƿo��9��x�i�\;:&5uFݙ��oo���! ���Gy�x(��Aj�`\r�g�bK�R�X%;��B�����=zgd��W��I� ����If�^��&����H�fw�xs��d�s�>8�����HOe>�^:)%!����0���l���IC�B�Þ�u�94*ʫɣ�ӌG�k�Z��i ,2"�o��&e���j�sw���ui�SM�9��T�^Yw8����F���n�V�xJw�\�#ia�!��֪**y�����c��GG����P�����{����k����{8'�`�I\RXXh�VO��K
Y���ZzZZ99���~L\��S�� Uhiie��=:��?Cy�~�4�Ӣ"Y�m��a=W�w�˥D%�Õt���3k�T|����_Y���ϊ��|����N��0���N�Ź>y��#��6��@L�f�s$!f��ݵ���/��U�s6gk�*Xs��i6��HyN�/�V�*?���|��J���s$o^�:�)�&б��kE������:y�]{��~��'=���\�Q|=��P*=�(ET�h9��z��/_A-��k�(Ű���MU��� +��srϮH�'�+Ԓ�'�|��w�����"���B��,����]IM-n`pp��i��p:����;��uuĎ|�a0�w;�'�@����V��#Ot����N~�:�co1�T ��v�y��6o#	��2�����Yh�>�HƤڸ��g��~ k�߭8���օ�h�y=ޥd襃��8q��@���*���)�gDuM�gǵu++4�GZ�f;�hhM�B]TX+����;�d\
�dʹk�6���nojv�R�v�O�S�?�3��QT�����h0''�|�dUUU�|���$A���ԁ(VTV^�;tu�iG޻y���F]\<HK[{@��6���+��;i0Ln��}�߆.��uv*�����~�
}-;;�j~~>p�/{��f�ߺ����\�بkee养
�[.�<ј=q�m���������/G�w%⭹�P��M�5Q�/l�X��#�J/�v���,=9R��ib��!�ŏ0�0�U��JY"�ԯW1y�d�>��r���~�A�}}� KQ����Y�'�Qf�*� ��`�U�LN{�i,TN�IkUH�2�����vzb�	&�D�ț�$'k囿u���M*��P�$�@�a-o�曌ʯ�:�̣�W�^�� 5���t�ӌsxuU������`+�����������ϕi�����џ>-;�_�U��"�/=0�]��(��HK6N�d��o��;�)AK�<��C?$�����J?���x��7�Y�9���`�7�2���k��T��:!���p!Q	I�U�h����~r��=ǵp�GJ���%��C��%TE�5�/S�=�|Z��e�s;Ҧ�Hr��̇-=�#�; ��T�=St;�Z5�w6���M�}ֻb/	p�=��1���FryA�eGr�b%�57`�������mq�����^�����h���I#ř�e�Z��J��YT���h�ݛ7�P܏�n���͚y��B����z	c��=r�z��	���������<a��'�;��?os�-Ey	��K>�o�L�K���K����}j����s����}jR�#��ӕ������7{��0!�|Y�����:,��8���!��0���$�)��'�2+7�V^��O�n��%If��� 3���,0j0TtlBƅ�c:ӷ}��?J�$��%���je����Plll(� ��:��.����:��������kЦ�u�U�k���-��ۓ�����C
 �Z��"ľn�O�s�~�^�2�pӼ
�O�L�ی�Ì�"����F�1�m9��洳�j��&�)��o����[3���D�[�gՒ�i��9|+�k�%�@l�OcM�j^۔n;����3 L��k��F"?U� �ί�@w���Zyv�L�蝖x��2�g`p��:�~(q@M=ë�Ǆ]��*�܅ׄ$S޾B��yC��o�`�)���`��Kr�ժ'��_�U"�ȅ�J{��;�����@��/%� "��X����߅~���1���C�hħ�{Tz��9p�ӳ��ԫ��v�E2�����^����O�E�T�1�g:�8P	:QQ��՝$�����χ���ᆒ휮�#����M|��4;�P��ql��� Jߊ�1����ŴK���Z��W�0�5�Q�A��U�YS��H/�(�?p,��8��;�c�95�u���4���0t����W��E3��Vc�1�Vw$�k>��6%�m�u�t�*@�h;�I襖ʮ�v��XdC�Y�� YlQRV7�W�Cw5u;9-�'�@u������+]F���T�]���.�g�/�9`{�][^.E�C'�֟n�`���eJ(x�5��my�K=��4�T���	G�k��Fi�QtX���nLttօ�7�q���s��ɼ�f��G�D�ꂅ��"��6~u/�忲�u~�|��������� ��'�5���K�F
�����F��S��)��5Yf�0�P�ȦQ[K�<���h��a��3���~@7�)hI�
j�DMq�����	�K#�(���^֖���R��{���I�Y���}K V��+7\��:cMe-��(�����p�N��Y~׈�d���$�E�a�*z0��SnFT���@¯܍J2��K-�O� Y,E�k�x���x&aK0���׃4Z|, �F���x#/��y�_.cʣ�:yc���zT.Y�����ʧ��+W�{��g?�Y�6�p����޺�%�X<]A察��gT�Q9���3�.��W=�6lI�<o��`�[qc����:��f�K\P�����#�S���ėYl�gF ��	nR��M���ɷ�m5Z�r�o��r�Ef�@�6�ֽ���Z{m��2r{�WV����ڊ��| "��o��e�K4#���6�V�˝�c�r����B&ԃ���vP�����@)�h�#���n�r� �p/��9��w����O.���Ύ�M��#/��r�d#�-����ΡB�L�}���D4� ����R ds�އ>�7Rz��03B���Z��U����3Sl���1�$ŊD<zhp{p&���\2���[�v�G*]�uϔZO��*}�Y�8NJ9H���ў��y
ľ�����{GE��S��k�~eL�̈���0�L��i�(��.�V�I��0���h���6� 	�����.V�⵭YܼR��=^�8`f�z;���\��N[���,��p�Ü����B�]�����2D�S_�E�?�6P/<npM��6/��a���zU0D`b�'vͦ`�Ѭ�3|~��U��T�������KM��C0��b��ݟ Ȁ�iU�+=�,l(�%�w�����d�Ms�rtl�4�Ga;i���#�R'�4yǉ��j�����ju@M~���H�֬��`�U�z�h�P��W#V��Wr����}�~"|��yA�-EŮj��S��oj����9�����i��M6d~K�6�g+��>}X��Ț�J�o�zw[���p�ЦHBP���68M�:�������dc0�뉳���;�7�f
���y�_3�6Z���;�xA�$�?�"W9�HB��廇��Zk��"�� �r"߅����AAK�vjQ:����?���/v�IJ�Q�����j���R��辕Pb�J�?X	�J�&&���k��q�6�3s��l���/�i�+«�.�{�x��b:��=���y�)[�J��n�%�@���Z��R�w�Ǯ7�7L_��I�+�9m*f��7nh�+Ι���d�Q��l��G�Fg./pE�����l?^f��$���M2���F��Gb�rIS�T��Z���� @y�{��mݐg^�h6���M�=�`����yI�u�h��n�4�l9��h�����V��x��ba��Z��:�V�f_�����c��p{�y�Z>�Z/���Uj�>�Q+=v?[�V}r\�@���"
�Ҵs?տ[$�,�	c��~�+��ٱ�|y�WD	������`����<��:)��f����?Y�>3�����S��9asuƄ�!j�s����`��m[�>$���ю��u/JV n|��p6?���j��0Q�8f_ߞT���2l��.�7�@9d�V\�>��g	�9! �-x�eo�Ւ��P��v�Ϥ�L��cu�����hH��x��7��J�Z�/�_�/��v��Kth�{�%�f�<�H8�4�zgů�H���T�3�J����I/7+@ 5� �b�t���y��4�p���R�pU�#����10xAt�pI��Ҧ� iB���F�x�$�n����H����&4��������Dg����E�f�l
.�:}��\yۖ0�F�e�>2�J_*5/FQ�@i�&�QX�[�沩��'�}5��U�I���![Gu{��������&��l�������V!�qu]c��A�3�\����LM�s��|�~毚��;װJ��LtT�����^ UQ
��Kv-N�kX�\����f�� CC���U�ݧ��=���tQ'IMr�P�;$��oE��!7��#�h4�kP!]�R�/��� �b�k���D	i�6^����9	u�r�ʜq2DLpz?�~% k���,��j�]�����utc�	.�x�[g�v�4z��w�ˬQ�t���5�t�$(FAk�׼����8�7���t���̘b魎�� ��,Op���IdmDtoO�9�����O�FJ��[��<I�T蜗�.b����5�S�Z3�C�C�>Zj$���H �Ԣ9��E�����O�J�K���ԭ�b9��=,-Y!R�v�V�*��yb�3#m��Pr~���E$�������
�ʗ0,Px�` ��q�S4���W����T���;;w��4Ζ�6)�vt��U�]"�W�S�U}���S8��t�K���GK���>! �?w�9��k�����*��7�k?T����kIv�NH��x���*i4���2�J��I���|4R�����SJ��k���v��nt�U][�g�07e��Z�U��^�x�J*2�+#֯;A�)&g֕��{$�@0���ô�Ù����{%
�hg��)�J��$!ܸ�V�n���NחKͳ,;7��Re��?u\6: �3���j.,��
����A��X�7)��#��g ��;v�p�3_&3n�`s��1�,�nn�D�K��|,��8X ��|r�8FY��aj���Hq�)�$ĺWmڳ�B��6�*�=�	؀�>�������9$7�X`.`1�5�Ux�Ԕ��M���o�:�}�2� v�R/T�r����۸g��h H+���zV������	���uk��F�^(����Y� �N4�?���=@<��l*�ɧq���4z��F,lu�&�������i�]� ��C&�F�pT]���W4s�zZ��׸��q��N�v�lú���F���ʅ�W<���<D족f��[t�҈z��1��W�����%�7�S^�]���y=Y�և�ZsX��gl�K�7�-�{��Lt�gZ5�E 򳍍����h��Ϡ-��L�:f��s"��_�<����Ll�����8�ׅ>=0�5��"U�r�@�7^���aC��(t�K*y�Q�x��.��N �����E���j�@j�N��5�)�M&�@J�M����<3m���~������bbh�q��dQl��J��厡8���%�)�<�I<HՏ��������$Y8ϱg��r-�/�(&�
��~�L��gS�O
*$�+���eAd�����gc�zݺeP5�����)G$!���~��M.5��&G�I�5��{n���{>�\E�G!���U�U
�&�`�AR��-JOd�a�jh�$T����ב��厙f��"�+M�a��.����� ��WK�/�&�3�?�l˴�KQ@��]�tzMI� Cg kX���$�8.g�؜�R���-����D)=%��H*�QQQ��-� ���*YKO�[E�N\߹ůF6b�A�7��豹<���E\���t�(���y�Y�)U��j4,�)Ԯ�݂'ʰf��ĐVy��a������GO1�SC�!F��"P�������~��î�����'�k�5���_8���V"�/��:��9	���7T+5�a�.��5�W�z���e�� X���:�K%S*��$7���"aAab�����<�%+��"���s���*���m�G�iw"?�,<Pj��~�W#X��g+�Hym�"��;�&;jl��F�(�\�ҥVw���
�乻�z���8�������dҺ��TW�y��I������=�7��-pA�a�� y|���
'���=�<�=��Ap��$?���������e�!N▜ץG��wb�T�z��35���	��c.s��^>�@3��avG�(_�:�(�J����H�ǋ"��3t����S䃀�����K��} �
̠�}?ac7j��Pw��/�t��1�u�Z�x�&�8�0	ƗF�/%������M��J�U��jñ�Q`��M����l���黷�vԬ��'�>;~g�h�˛:~?me|�˴���̞�لN������&��{����K-�p������q��E`�Mє�ab/ ���0k&���.���s�	�9ТK�ȍ�� �N��v�nQ(ȞB����S1꿒�yAH�/���N�!�C�U��E˃�`�>�Ai`ńDx���<J�/�ږ�^1�f�<)i�l��`���J�o3�T��j*�0�S�z����hv��)G>U�/OK�C��$4�ǂT����9e;|G�sY�b�MY�N��"�G�eY��@�#?�����3�╲�鉍��p>@;�>�?e�y�A(� 6�hr����)9z܌�V����c9�����R;W����i���p�@C����I4�b-;cW��M>_�y@c�g�H�x�b�4oP��#ߎ�����{��Cf����Փ��?»`܎M"-G@���kT�ƌ�"��� 6���K"��ι�����lKQ�$M��������������L�Z�
g�c��1bC�Xڈ�ΘB�:S-��"�}���y� X@K����y$����SX��@�ēu�A�X�	Z�B��)�\���?��l��S�������3e_����Ú_mx����H)]d�T.s��D4B��ɗc9��< 6)��?�,]�ZP��l�
�y߸�m����A�� ̀��Gr0�a5���#[���4�?����qH��I��L�-#��Z%�a2�w\�%��*ۊ_{�~�TQ�h���pDa{ �H�U�R L� ������꿲�jS�uxq�:�ul�3n\ž����Ti�
^�d�4���&��밼'e?齸lK��2��CL�׭��dڦp� )IɁ��������Z3PK����D�5��Ŧ{ip��7��S|Vd�0 ���'EPa�<�e��b�����A�0�Q�Z�������҇�r�`���������N�vf�6U!2��7Y����DJ[?�ww�2� �{#��)K׼V�&�o�0�S��D�g�Z�nc֩4�b����~N���_�J�~����ߔ��V���dZ�g���x��Af�Ў�;Ku�j���"���ګ�2��̳6g�Y4���S�P��s�0��Ŕ������WLH�`Jnʁè����#棯�`C�W�6Z�Εgп
����1�sЗ�%��In�y[�^ǹU��O��P���FJO�R�[��O~�U���p�A���P����#F�:�`��+5O��f��g�᧑I�i��� �cIu��ۢ��W�/�ð�c�.[]6b����>، r���*�l�S	�]�
�4�;����]S]��G�{�b�ޗk�O�	��>'`��+�L�T�d�
,&�&����`�q%����I�`�eY��V�������Sq8��t�n��wu�J�B6���Ө|+	:+'�}��o9C/�{�U��cA �]2e�!���d�宝�_���lIU)��ܓn�4�>��/k%yr�,�I ԍ]U�J��.OJ��O����7�2;$�����,�R���\c���{Ū�~�MH �+y^)���h��8�6.}�'�ݼ�,�����f�i�����#��G����;�Hʦ�6����B��w�{8�q�Z+�(W�ڷ,�ð}Gas��t���(��
6D+o�㳢Ξ�-5p��o	�#� mܔX�.z�6Gh}Ʃ?���F�߽ٶ_�aن��O)�W���%�̈́���M�H�.I�'Oa��ɭ���߃)�q�֣�8�ttϧ_ ��R�3��C ���+b���zj���u/�A@���џ�y���ҡ�u��>�,!��X�b0��>j�q>�����';�q��{� �a�
L���W����D+ye��J�^�%�&dԲ����pE4R�#�l��L^�FE��	C��vg��O	����o�(���P������p������ �N�S���w�랇�)B����{�,����}[�4Ö>��y�]>��1�����=��K۟qd�Y2��R���i&㤅!���yǻj�ŏ5Mp͆�D��Ͽu�|���sL�Lβ*-����΃l����!)P?����<�O�kn���3>xL�)W�ɖy%-B�0�	��wF�H���2�3�.'�=���q@ގ�d��l���[${����h3G =Y�a����0�\�`�d��e����wMy[���(��k>�(r�|�J9&�����k%���S���/�]t/N�
�����ax$��X�[b/�E@x��q��y~�x���)k~l��K�H�j�IXϫ!k�Ay��_�b#R�B����嬡3'�`Δ$rO��� n	2�Սf��T7|Rp_�^�ț9�j����e	�)1�d�|���m� f�������7gI�K6��%��jC[&�|��[!/q�� �JC��+�M��mu����+��&���أG	��Yz����fɏQb����.|�M̬��}��6�R�͖�uڸ5��8�Xed��l�UKRҲ#�$�@� �<��h�fS;<�����	
^�j��L�Z.Br����#�U��;����5�XT�ޛP�)r�	��y�;qC0��e��̪6_G���[G�ǀ���Ӽ��VJv���U�s�j�^N�h~��u �V��{�>E�؞�{@]�g
�2�^���bN5��q)A��� �v(n�(�U���wO�I�sɸ',h�<_Yy9�e�^�`��h��r�.5k�g'!��i���#�xƈau����w���]#^�mI�9�Ȓ�}lZQ>�B�tu����H��H�_݇��ә�L��x����s��!$���X�|݆�Q��^�q�&��9QD���]0/��ff�<N��D�Y%� �'�W(2�#��^�b�>�����fh���ȗr�Z��ޓ�nu=k�߫����s����siP��|�/�˥��9���G�RȚ0���ѾL �s��=���eS����ۿ���>��|�D]�d+cy232�2�6�BV�^�Ql�[L���X�>N�C\*IV�<�@�_Gn�$�\�Ǥ������� �o�٧�����1������I�x�
�t�k��`ro�L[ʩR��C�)3��Su3zp6n�@G��$H)��U6x該Y:,gR���W���`�����@��G����).�����A$Qq1φ�J���B�A�keV��� �a��+���h4��Ie��9j��j��[r�}u����\+�D�x���>qFnO�J	@�s=�� ��x|[RNI-gu����wcw<~�iJ��Y4�?�4�`��dV<N���Ɗ�pw��&��Q-�y��i�x���q���������G%ݛd�fO��Z��zi9�z`�Wo���� �(�� �W�4�V��;���T���[D�����AAa��{��{���f�]K��g��~���w�K�L�5����k��g9* ..�Q-�즞'o ��2��>0�F5'��9��Y�.���������]��7_����?Xv�ށ��`hY�_��{�?�J�,���rL���y&t��s
�3��j��I�\iu��B�����2��Z9bBuk��G}3�L�a	=�Lـ���G�p���jo\��$|�>H�� o爩��� �����sH=T%��X��כ�w��z�01�>���{��<�j��!k�Lc?L1�.L�ʝ�J�)�<���zG�#�b��,{T �ssG���#�`^�sz��ҭ���{��-%�B���z�^3s��w/UzWpp�Ԇ����]�BpH���A�3q7���}S,E����q/zR���Qb�;Y����%oI���C����փǎI\"��j�{Tn�q�@	�ͳ��\K�m�T5�D'���Y���C�0���h��cU���^TF��i�[M��x&���a�����Ý�>�׬X�:nH�N�瞎����M��Q.����KV�{PdŃ/Ӹ	�5T��nߛ
��d#w�����������u�P�:@��b�6C^�-����;��?SJ9��_��M$�	1�5O«Ȝ!�I��ř�"w��6 �����6�>���*� X�,�hs%�� U�$��$���E] P:Ճ��T�FZ��+����4�,���>*�a�s���!4e�}'��ԿJ��Q`�A*�y>�6���%��7�"_@-�:�cJ
��f���1)�Y
#��������>��<�+3{y�o;�2>&����i���ս=
P`�-�3�qh�P� �i�R�V���Ǎ�:��wD��v�9��2���#wd���ڒ=���h&�b��Ёg�=�L�k'O��Z�)�� K�Y�dWxI�M!$_��x���c̔��_��Kc2�a���lˡ�?�ڒbԂ�u3\�X�M�j&[����+��S��ގl{�����u��骧��!N�-㷙���sN�{e��� �ڢ��7�dV��/Y����!'G �=��m?��V�<�J��Ӵ
<m���ω=�������!Eg�:v->}O�u��	2`�����ďI�5��u\�U���"���H��2�7[�A9�:�U���+�|�u�6�cVmb��o'j؞;�K��5����:S��ȃ�/�����^լ-�~z[Y�k�I��gV��} �{��8O� ��`?;�cI�9G1�����/&?�`�l4���W��f�-)��ZMf��^e�!�y�58DC�'q^S'��T\v3�0���B�Z�k;���x�y5�韼�DY}�V��2�j|�+�?�Z�:փ�?& �	@s��s����Ȍ Ypg ���,�f-$1aXaWs��1>�݄�$�-�����Lk9��r] |�#�f��sM�:gUo;\�
��3�0��������5�kҿœ8�� ��A���Mc��e'KdOFB�/���s�U��Ђ�v��j�	��ǾS;��?&��xཀྵ���#�x��[W���\�r��#���~a����贑gl�
��~#���
���r]�[Pt2b��57�F�W�fs��t��X������FR=~�n9rc��N�0��Z��]]/��S믤�u���㷭�jmltl{$��śH�m�����8�9g̃.P�N��>�ܓ3O� P��F��x� Ӣ뛐\Zrq�K����]^�lDP�ڹܨ���Y�Q��I��3lh6/��׼��	*��SV�%���S���t��1ۥoa����Izp#��^���M�RHV�l§S��hHxc�ໟW^v;�0��D?y�Q��m6�2�kf�Q��{$�/�!��0��(��Z�k?�m��;�p�V�=�x����% E�g�DP�S�fo$�)���b�}܀�ۨ��u����Y���x�Zj�4uAj�������d���Y��#'�6h�,�cݜ���$DU�/݁�>F�����R�q�����][��KW��s�5����$�VI���Уm[i���
XCa�/��U�mRL�&%�^�N��'�(;��>߅�#�d���j��v��_랻ל��P\zBjx%��=��a̹�;n
2�x��/t�A�Ң��z��̿}� �� �'r[ȸ"-��j��%+�TW�6B�׌�an�W�ٗ���'�x����e��M�/�p�N2u�&���) �3q�Z�!-/v��b9q)nxXW���Վ�s��X� ���������dT�Y��?��� ��¢��5�!�R����M�J�X>�
 �x=�Z;c�f�䍙�j��-��
�E3��Bm����S�!����ͧj��߰��.�zj�'�V���z{�#^&�b��d�>qȋ��㊩��L�ΛS>]�}�F�	� X�u��i�x*���VL��������-�`���4Ot�*.S�޹�,�@�eL���V��Q���v`����E���o��7)���!.�n`�� �5�Vw/Tb��m%�����S��u6{�
��k��2�~_鄏U�x�C��=��C������D3.Y����|q�p����E$y7?�C�d�F��W�����b�?��E9�BG�l�wJ|:M�����yT��[6̫C=�o޶,�����D��s���w.L��l Owٓ�Q�`��V�7E�}��_�DO�|��j��$JJ�Bh"��_?B�����؍��[+)���KR�60e�ڙ1r��)a������⧳���R�b�˸r�3�������Qm��CO
 �rk���F{�1�V�M]_go:����������������� 2l��Hy�e�\�9���|��H�X|!c�<kV��VN<��B�p�5��MpQC�e-ҽI]� C��.70 ���_���i?+6�����-���<��j�־�\G�;���Z'xgF�Ԣ��IK�����[}���F��ڐ".����r�A졉���h�}bYX�w���p�p]f��w$[}����1	��vWߣ��;ր*��k��+�����d(�w���V��ئ�X��Uq��i��8)b�}k�BY�L"��@38��0�3t(9��1<.e�u��ʛ�0��T^V�J��,I���v�����S��H����H
k��޵D�k�#Eǐ�Do8!<p�ũ���ٵT��/I,s#_&s���<����I�.l1��� �j/Cq�ֈ���-�/t�I��?�Xm/-^릭r�Koٮ���-C��W)�)�6�H�_l���hnq�=||���Ǘ�2S����,�e�J��-p���O����\��8US��Sv�_;���O,(^Z=i�=�}��b�����".d�jt�٪�[� ��	���������y����z�J��\���'Sa������;��\7��Ȱ_%!�t�w�B���O4SM�N�� �\��9��W�HV���OM���K�\��a��ė���x��pʆ![�%�:����?d����1< T��T4��3�)ۡn�P���>5�|^�p��@⬨�4������4�3�2�~��_�˯ztn��b�n�X�F��g�����K�<�8e�F򵓚<��b��鸿��*��9��5���+���M�L���l���ݖG��G,�h�������7��#��Pw;Q9��
:Z(k��ͻ()z��c�y���䝩�T� 7y,�_x�|J��קѺ�H�ݸ����6)	����hi�2b	�,,��Fԭ�NWx�^IwV�&����*��I�֐��V��DE�����ǒ�O�^�ޭ��i���Vɗ���L_��j��oy��׌�8�����k�K���JJЙuc�j� 9Q�O�V��0B��x,����lt(��j4�$���B@]�JԞ�v���y^�EW#S[�.uW�j�%\����p��\l՚/2.|��V�wf=֚� �eG��Aǖ����6�1x��ML��u%*Ѷ�)geVe�eQ�XF�%r0��K���zi��a7~��Ϫ����6̞���w� i�Frw�L~���(e�q�7|n_��[���ɡ���e���a�Hš��,]�Æpe��kjVT ��ӈ�Ǵ�Jd���x��|֊��uUuF�v�3���c���^N�Io��S3����=�G�����C� �����t������-�X�a�"�����B�������[<g˔F�Z�%�"��/	W�e��<�g=���O���)�˗bG��DL7V�i���G8���3�h&�����}*ɞӧs�]�ItA���,�����he�3~�r�>7����Z7��.o��Pm��j��UҪ�*Zp����O�Ӿ���y�v��cI64H�g�e`����F�LC�Փ
Êн"_]�W���I�j��4��j5(���}��S{��̙Tsl�����r�$�C=���+4�,RF%~�g����:,�uR�MHjҖL$�ڐOV��G�Z�76J���-�l�[e�c�l��f�j�����5ˉ\�[4<���y�t]��Ë5!�$r��ߥqw�
$��щ��]� �!y&�����Xl����V�B�ن�����;�B��\����yA����i��v�T��xGz�:�$@�(3�,���GV>w�FXk��� �瑮Y�-ѻ�B����ڶ�J���]F��k[��K��a%�t܍�B��D��,4"�r5��K�G�:k�P�cU������X:.�;O�ט
ڒ���a�����~<fbA��X[�w4��`���&Q�O���l����H.g��^5��?p�w=)��vU������}��*]t���_O�I����d7���VK�q��	G&�}�����eJ�3N�x[�Ζ�A�<fe��R�2���r�5�s�����d�-��DI�T6P袣JYբ��fIz�����r�rz(?�wE�������C�W v����l�W� �n��M&
����҅���Y%��>9�)��㮪�wx;g����ȷ��}�����a��M���ಊq/�����8���o�ļ�g��q5������^W�i�T�̆ њ*Y�Mp�?�x�aXb�3�ho:ju�=�C�ʲ}߬k�e�"7g��t�C�3�4��'Μ�)���Mo�鴡��7�@٭��u������l�f�C���mr��ӥeÚ���w&+��k;�7�yM6fn�O�_�4�i�/��_�1G����/�@w�xa�7���)�u��f��|G��y�%U�np�L�k+���~/ؿ���=3�8.;����+qI��a	ʻ��KQ��$��Z�1YM��}��×N2�u5O�L�_�ļ�J�w����-_�ua��$�\l(+�LT������+�cmQ�"�M0��ђ�1)��h;7�o���$�?�@�E@�4)����?	Ku�ϖ��Q��;�Z\ibW���sV{�)�C��`�X��M\	���zM���r^`��;Pkȴ'�r#W���).������5�'�T��\�7_��Wh�J7OGdK�Y�ȮᕨY��X9����	I�Z�aiSF�Rړ���]��s�F�&��B#t������k+xj�A\(l��>�JEe>K�w�DQ�����M�yo�������/Lk�֌���?����ؑM�Ԙ:]sӏۖ��Y�ܽN�E�����C���]�����G����\�
7�MǇ��,�8�ȟa���a�ݬrt�j�rJ�/�8)M5����C�=V�0�(��X���ߞ�.U"/V��tV�C��=��H׊�0�N"Bdsja0�+ETX���.�Q5i��°�v�ˋ��ߒSe_�\�g]Y妛M93��9��់`�B1Ӎ/])��|�+LT)�m����E(F�X�<f�B�c��KB����(���n>,!Ry��P�
�
dH���f�i�~R����d9X��A!'��*vR&д(&�Q��U�to*D�<+�<�W���)%�h%,����ܻ��}F#;���Ĥ� 	Uc���Y��Q�����@��Zv����usb���cw�b5�PW�Tz]X@#� ���r����T=��Z�,��j�9MF�}�+�xe��ӵc��/J��\�QW/�2_�l�c����U�+jXh �i�ݵ�����%l�vW5VN�zg��	���1��N6�? �
����P��dǲ���c�62���Q�F�X]B�|�F�G\-W�5�`�V��a5X�p�p'J�~�*�bإX�֔M	���{*D�-�Lߗ���5���i6��e������g��q��0%ɡ#\�����ٓj���F�Zl���U��f (y3�2'��Պ����_6\}�#�Nѡ�ϙy�F	Q4.t�Ӧ��Fp����c_bɗ��3K��k�ZЂ��o@�
s��^ۖb����e�K��H�0(��;�8������T�u�#/��޾HS��[�f���0��'բ\̓Sǿ:��ػ�M[��X/�O�Y}d�ٓ~��̕y?���C�bV�@>x�ι ���%��c�z�~A�>>O���Қ1�.忒�o����P}��Jl�{}ե�jp-����D Sx�C����>�t�U��`���z�Z�_�+��� �󪳩Be4��\��ol�|Oʞ�ܧz���/#f����K58��!Z��^ᤑ������~��h���K�@��υ���!�������˧��E$&}��FM��y�\�x3jnݲf~ej�V汀t-��>�}����P��M�77�S_7}�3* �ؕ�����7�q���v�/��H��%~7���ԅ�90�.n�:c�ds	VAM�L>Ɓ��Ŵ3����sunof}x=��J���1I)����+l0���"�O�P��/.�$�^5����<� ��ȳ���`��Ԧ./6��eL���i����ơ��.͔8�f!���x�Y�a�n�>�SFy�����N�������L�|��&��'���c_�6 �&�k1�pև���a�KⒶ��+�kr 8�*9t$�BP��^"@�)<�{>�������Q@Gɗ/�D����a�$ �y�Bs�A����ᯟ�-K�}&_E���������Hχ	_�n�q�'�B���B������濾]�\S���7v��(6,o�H-X�{�	t���͵�ؔ�t���d&���c�A� Jiͨ�ɗ*^�>��[yI1���4�D E'�����ڔ2Ta+�R�L���Kf����̣�4�1����nh?���a	\wF,v���8Bd�ˁq�y~׋�/ {�7�M!M�	,lJ�Ǽq����s��H�g����C�yx}1tMS@�.��!U��/W�ڃ"SR+hqh^;���/����ӕP�5GgE=���Ի`ݒ��v��t��"�c"�51OB�&`��/������йu����L�rxWΑ��/CgӄC����MX��i�%�?Xw��xj�w�j�t�-n��.	̒+/�Q.�'瑌E����o�
�Yq#�B��xy~�0�� yn�g΀�PQ���X�{��L7XT]R�e� ]:�E� ���ڞ�&�+���H3kVX����/�
��iBO �oS>&��><�rL%g�-�{�݄m
�n�7ۼ�4VK|&v�W������3��;0}����V�F��^����ӛ��i���7}0F0d�=_E&@��7ł�,]�]��lH��\Ј��(b��b��f�+��;w�Z��J�D��i�m$=��s̑Q�C���yh�}N��'�����c���C� | �	eA�����ε���tǖ���"�ڴ{]��V}��O#>Ȉ A*��x�U\Q�q���+������J�a�-����nғXuZf���스1Cmxh9�����jL@*�)�����&�(o^���5��4�U�:��DKu�g��`3{�Hf���q ~��B����|��P��*�rW��R�S>��O�k?���D�1~�v�������<!;�f�9x�^�nG��c��)�C�Q��e�P���|����T ?��m�h��$�|��s�ϒVkމ4�,�]�Eс_2=߷B�~뫄N熫~�c��*Jv;6E�;�Q��9ru�c�.i��DG�>�oJ�_	V�FҚ�3y �:�p�>�-��G�80X��)�>�\}}��r����jw�|����K ��7:'B�4�N��0��b���C��2�Es_$��Ze�
cO�f�:�;���Nl;9?K�1���Fs�l��>V-�!����L�a��,@,�vN���ɝ-�N���mcGF�\��r*X���n�[�<F�'�%-P�9��[[��[�@5Y��d�Ł]f���>ǵ���оB�����؇�%F^�t�&�)1]ܐM�*4Rw���X��t���S���S�#����?�o
����{����^��k���`�m-'�d��_
md�`RJ1�.<�<^���R@�Vm�vБ�1�!�F�#���M���uYN �E�����	����tj_1�:f�KS��iW�Α����_�BXN���A^1)+�ޅ-�?d��<����i�2T���)اί�����6��yR��7��3Z
�9�	�5x9i�J�8.@�d�L���|rʐ%�G����O��iZ���^a�0i�:|ްt��/*�;c��[�"tT ���/J�����Y�@H���+=�<ŨMm�@75aͅ��
�i
��M.`�SjSٚ�q��8�n����Zz����y�Ou�t�H��'�&�B��a���d%��A�5 E򿩿	1�N�Q]��ҕ�dͲ��<���{FV����22<("�\�hH��_�ȋ�L���.���,撿=d;�.U�&N�I�	��R���eTw������D��M�,���w��ĵp��[���/� ��-@Ҝ,���(d�r��>���mc;Kv�Q��3=�J�)@B�h6>��C�/l�a�OC�jpv_�J�A���?S��C�YC�:JP@���T;���2�~����s�0�S�+J�����֥�.wVU)�q�=���7w�1�Ώ7[��1a�Γ׎=a�<���g��!�V3k�c[��c�7�Y�;Ĩʦ�偩%̏�,����$���ԇ^FQ�$)yV���e�����g.��\h�V�߾���d�KS�.�i��w �X�lb!U�R�1l#��ݺQ�ݬ���=%����s�F��ܣ����s�F�P˔�k��=֬��ϭ6�G��4
�h��5��B���� ߔ.w�!�[X���MN�S���iG:�I�p��`�cn�݂$g0
���������5�$���E�$�&���D%��К拿s�& w���5*��j�-�K��J����G�RҒx���O���H�!$X�I��t��h/����}���k�fژ����)����Cc�i²���� �߯f�!ȵ���ݱ����]����Gj%�5:�ix�������gC����6.�dZ��~�x�2E.�T,��Uep���/7oH�!�tf��T9z�N�=/.L-���F��|x�he�i�ӎ�T��\rK��L�狳�5�M_ą�^$ؓ�.Gy���=/�W.,������w�������b�K�:�Ug&k�ok�Xfn�Y(��Ӳa����
��+c�X��:�6:w���p�E�b̢��w��Lŷq-fZ�vn�>J@��2@}�	�4m�Η�@�����;oD)�1Ԏ�O�P��?�ک�5Zd`�Y�-�K��������*a)RA١������:�o��=�O�3n��5�&�vh�ٕ<��-o��G#L��8 %sљT�Ցu*���z��O��+��(�r��Vq%�i��#p��f�_4�wn��� ��p�c�c&��:� AP( K9p�����a]�	�1a9#�ze&s�
!S��}��eP�����4T\\�jťƤ�>�Ǳ�b�,/-Hp@Z*�$�;�m$�����՗����j5�};�������u�F���[��4�lz�O��e�c����	�D � �^�l���jG?���!��+ݼ�z�R4���|$E*��@��W$U5*|󿭺�Ӣ�V��;/�NN��y")P�����dCԄ�*bF�����j��,-���8_�������^Yf�O����!��1�rX.�xo��'(Z��Bi��Z;�G"'޵R㺋&|��m,�I|QO�f2i(}쏕b<�oy_� ��@���i/��IPL�̥r��x%�)��k��U��R�]Ԝ��i4���b�e�@�ha(�}P%���CH,�\����J*v�.�
����4�j��Ƽ���4۳ϳWͨ�UĨ)Y��r�[W����0p�*���*��6be���@k��Ƌ��G��t��(8s�kզN6ן	��rW���jX�j������@�r+�^�qu��$y�����������i�UNm�GN�ú�E����F�ԕ�ǦC�T�v	Y�	�}�ݢ�і=�7F��?t���l�pk�g��<F��]O���v��> �N���@�-��|,T���:Ƀ-�4��w��a���/�v���J5����y�Lg���_?�,_d�d�VP�ü����ĮM-��LW!E����)B��#�Up�M�i9t����lI,-��k��T��t\92�g	0�i��*�dÃ�-ZU������FW{�;�%sX9j�腺����YR�>	o��m�9ɬ���E`�4e���(�x��%地`���G�!	\T9yv����!?�M]�������\{f�*Yj1�Ez���r���h[��&�$^��fG۱�y�Q���ǫ���xh��U1����X�Α�wm���7	�w,���ܧN�|E��Gy�s�2j�V6���/��kk��t�;C�6S�]���3G뺼i՝�T�j�.)����0�5�|B����Q)��y��V۫��H��ȾUZh+{]Z�Hǣ�T�R�\F<��t�I��M�흥��Y�;��XY�5��ۮ������yq��c���ZkX�K��<�5�]�n��� �$�`�G���Q	'�ms�=���H�S��*��p�!���c �Q��h��j���f���y�U�ֱ�;C��ڍm���V��jW�+����'ᵛL9�ڧQ���ŀpY?��[��
�o>>��un��7�c��>�]2/���LǗ��re��R�iRD��uk&���%��qY�s�&Y�����������%�<�����$�T��XM���l ��ګ	vړ⺸o���{T5�\.�6g�-�A�_��|��B� ش�h�'�Y��O�� SZƨ�@�M��f-.��[W����O���a�����2_F)�~}�����ܹĺ�b Yv������k�0���r��c;�vm�$��)������hn:E���xT�y� e,��?�[W�H��:M'����a�B������SH�{�.s�fEީ�IA�<�`z����ax��d\��%m[�KA_��m �pQ�>ƺ䓈H�D�:���R�|k�j)���YKk�ݨ�Z�Z F�+QpfGX��7�X�6v�9o�hP汍W�Vx&^�%}�f��-�<��>p���B.��?}pQ (B��kP��m^����B��x��!0�ѫ6�x��_�h�w��L��f����a<Jfl�~���w��ٲ@�1��z�!A��A��O�y��!��v(�"<�� �����c�̗�b�(��	:�c����}4��:u�Vĭ{O�%.PW�o����Xb
$:8t9,r5�;�L���P?��H��c��Ee��{c���T����"ڜq�,����敐���s�0�Bn����)��'����2�gk��>oV����B6��"?K�8�7�AY���Cא���S�nG�඘���V���^ѷXϴ��\Oq��RSb6��X���������)\�
}�Έ��r�����X1��/�����G��4w5�v8���k̜�`婛�Ƥ�����2��⼹$t1;�B8)T᪷�]��6gE|F�� ͂���G�k �$D�TE���X�N���#�ׅ������F�C���_��,_��2zi�#�Sh�?)����a�&b���Z��sU�ێ�a�d6G��0�|��J8	hG��Pu.<Џ~Q���"�u��TpW�L�x��Ȃ
�i�`�-8/�}s>_�^��U�i	��6*uNYi�-����\����w+�Yw PT\�������|���]��l�߅�hi�&�Ŧ;�ݟ3�\\�3�{W��C���m�ѩ�wD���"_P�)l��T?/uT	�"Bvj��"V��pv���ts�vk�#��C�����b��ܹ��z�����܄m��яg1�?#Lrd����Q>�Ypw�r6'�5D��w��Җ����
�,�;i���O�3qԤZ�ᓦZ#�C�q������:����/�n������Ғ-��7"��� ��t�D�q3�o���	���[uoP�]��E~�����z5ռ٭g嶓(��k�^&%��VG;i��p�8�ؿ�k#M���N%���㦲�'� J2�Xa��Hn��[V���J��搣*�����!�\��`\���:Y����5�
�����t#�%��J@e��r��d��}���]7���YiU�	d+��0i1V���\����s*��5�O�?��p�B�\۴q�jWV�����j��3���?�սC�o�_����'�[��؉$�ܖb!#�����顰^�<-L�s�Nʎm��m��ݵ�T��ǲ�''�;g�4x�ۡ�L�l�"�:@�J����6�N��@��P�������<O�Bk��gm�tm�a�Kn�f�m���r���>}GVC�}�JD�f�d�P��$g��\����+o#��<x\?0���|6�vј���ުަmb�$�)Γ���Z�vJ����]�Y� ^v�,�2R����q�"k�E���I��P���>����0����9[�lH|z-�
̬��@^�	��r=���K�Ŝ%3��\���*����@���+6=br�3�W�k��%�������L��`ak2ׄ��!�	�-���lHQ<?�Ɋ�o6��� p@Gu���_��B������#�W�U�:�YG�خ}���|2km6u~ۛ��ܟrR6�N6��SL�!�r��t�8�AN�����=�g�8��h� �ɾc����9
)�C��§��l���'��ە����PÃqV�o�E����ݧ}	$�&�>���o�<��]�dP�V�!Q�!`���*�Y�l�uɀ�I�uq�nn����5���w�K��I˨C�]?��`�%�G�6����!D�E��t^�z_�=Vɘ�m�3��g&�3�f���������������C��Sg���t���0��1}QG��0c��XX���d��� ��Ѣm_��ˑ����'�u�i���&`~��=D�?���涋�� y��ohgQ,ԡ��g��������}
m<~��.R�n�Ԓܒ�n�2�6�_��6�m�����h��X���QG��}&v{�^7���浓�T�L��K.�VL�ݹ����
E�!��k}�s��o�b�Xb��	~�ɨqk�b1ц��7�ɓ"^e��H��ƶ1�-�Ҥ�SE�a����< �%�LW�Qk1�D±XRP�{Y2�����~E����D(I`oi�����)]"���Z^c����_nF�����r������/������T��v�#�aʁ��ҷ��UwsG'��eT���<g�at�.��5���HxN���,L�d�
*�� �.v5�>����K֛I����m�R��
 �72��l�D��	6vSGe�f9����W�*S1�X��Z���q�oV.V˖�?�&�q��b��+:^��Q9�(D�[���Ϳ�r�;,e��%vh����RM�^�i����l�:��*�0"q�RX�	�zp�N?d0�e&mxG�a�۬��>�o�#�F��a�q�CZ6��t�h�m<�︋�d%_���&P���}���k�.�s�_A��?���ݱI�"N���'�?�	�tx1)+;)k33='�UG=�܆�c	����pnx !4�F���bg�Y�/�V�6�U��u�?7��lcG�*O(!k.5&�q�����9�\ZLI��N&�.�	�89�L6V>�˖���䨩(X�H�C���O���rɣkWd�X��i+M�K��N�f����ʩ�hw~Vo�kh<�(�����'s�GMea�nP�.^[[�$i�o�Ts�������.��m���_�Q�&��z|h@�%�c�v����0�5>��s=�!�⹡X*�$Ӡ���Q���e�v:������۱���BO��|>�~/���1�������(5{��g�l�_l���?�WB�n���9�5Pe�C�ǒ�}%���=��"C�(UzU[!�C��g\�t���f�d>oж+��Œ��&sl��:
{�]�,�W��f{�V=I`��3�` �l���-���j���h�2l�n76�ߧ��:p���d�υ�s6�q�Y��p��<�g䚕鵼7{|���MX@f��6��qr�����`�|?���>����Ә�?�O���)�E�"[��Dɧ�<�$�\��>� ��"�J9���.�o��)oZ���;PyЄ�F�7Zn~s���>��;��8Yf���;��uO��}o� 
&�q�ޑi�kO"�� |�SR�M��i;k/u9�.Z�
�+S���� ����r���~}��2Ci0���
����e��f��Nq$�pf�$�J�!ҳ\N�6���Ra�5���|S�U$�~�� 1�C)�����2|��]�%���R9SU���?ơ����lxr\�7�d��]/��_�����38�6*?6��P���8�xE�f�8w	��Rt_��\O�o�`H��x%D�b�p��7H�}V���R�p�C�r?-��[��.p�M?�)�Kr���d.[#5RnLԃ-v��8l��?\v�}Ab��B��k�כF����wG�"���4�TU(d�]&÷Q��WV> �,AT�;?{����\#3T������*nGa�4�L��UĚ8��E��bu��dՕ�4q}��*�W����[��
w�3$9I Pw*l3&$Db�д��YQ������PUM'M�	>�d�T��N������ڍ家�m�vZU|��h��k��������s6�@�0�v�k�(�� y�c����/X��mS�T`��O����~�כX�K��H<��H��i�*��i�(�i����M��'UnJv���#w e�{�Y�5�|j�����n�2��efL��ܟ_�]��o��N�q��H��u��IuH�_��|�݁�*�1n��iI��q!hu��ct��W�l[�s`��������[�гJ�=\�4�T�-AA�G�I`�[�����~�2`�"��N	�F5+b#`]>`�+��(^4;�Y�d���b��ee�v/'�3n�gms5���B����l����qN��lﯲ\��wUsu��@�K���	}9�Q���(�X���1�s�3�޾:����,㟿}Q�XE�w�^i�������6[���<�6�|sl��UCn�+t�����y�(w͙ctP����������?�F�Fw�"��Ϩ�?� %�
FWs���z��Y��[��:��/ʵf<8�ϱaկ!C�h>�4��T����*��N�1�U�J�c%�8T*w&b?~�����?�@݂O|�r�V��h�qNO�x���v�����朰}\�J)��Pܥ�e��Y�I��|�����B�i�x"d�z�w�gb�QN���q�5�4D����	�M�um>��~gTQ$ӆ�L�K }�,�=�5̏�UM�~�;�7ͳH�[2���U�S�3�}gݒre?�O+����aH2��-E���@¿y?_e!����~$,��5);�7w'�4X�\��:�t�S��(}���"e;I�,�t����咵�/��XzU.y�n:8�V�6�۳��V)0�6���K\�μ�H<��P��#A�PT��v�0�����s��c�^�@����_j��{��{��P��}�<���x�ap�>�ff�ӏA��4��Eë9=��;��Z�@��a�@���U����/xBy�T�f�������	? ���H.�_�u�[Z�ǜ�'\�V��:o)�WEW��uD�wi����΍&͂�v�ro�bP�G�)`�Ԯj|kc��svDu�u�<E��K5'lE�OՓ�T�����F�g��@�(�p��/�C����ԏ���]�Ӳ�	e����g�i�2p�|�"Vᓂ^��t���b�]��D�)1w�h�U?;�?�Y��VJ$`�v��}�U�����7WUe�dm�R�%�秂T��w�ԙ!�z�1or�����-��0�lC� 9�UW�|6��ǚ��@��DF��Y4��6���WQ����>0k^�5hK.J�>jw�]B�Nю�>�f?���z����<zG�5�F��M���4�߈}�_���ztz5~���+��CF��� e\z0�}�\�m\��e,��$9̏�s��_ۍ�h���=y-7�h߶��9w.��d�f��v,g�����;>����;��w~@�|���eo��+�sgq�9���*��&K${���e�4��C��������[�~�s�l�h�1����i6�#�o�:����.�{!�����`�[�!��xc�	�>��׳�	T+2}�1i<j>[z>�(I,������<
����Z�����79˟-��pw���/�p5_���ӆ�-���P�}�_k��Q��j5xЍ_"��T�1�T�b����*ϑhX�"����W-��{�ݿ�%Z� �41��;A�� �Pa[1Mw�DN��Ơ��i:�ru�%�}��<�a��<홇	���.̔���s%���������P� �My�����3�0�,��&s>��s�D�y�[��o V�����0���]����O��H��
��~gwf���4�dB�7�zq���@6�CY��]�#	{J���Yު��gO�k���;��O��{P�_	yj�E�ݩ8iT����{4���y����whg�XAR�s��s�@�˧�ssC��:���k��āF|�������
�(CT��HC_J����缇�^��k� ��;�7�o[,n�詘�ǈt?�aq�n"V�74C��*m`���a�������̰���0�m��9�q��?��;��r��'��y8j�X$^��@��b�9*��k.�f�3,��۵+>>SH���_l Rt�9w\�%rl�p�ju���Q�Y����g��j×�i����Y����p�ƴ[�Y1w����v1um.�pI���Eԫ�2�o��q�E3ī��D   5>���rl ��brY����Kt����ϥ���(U_R�rc��w�;<	e`�#�����3�E>����5�*�M6i�n���t�d����O�Nq�غ�@��3�&.��U�6��3�����x�.���� 9�E�^|Y�9^�>׺:�_�#��&b:˥����S�QByu�C�R�*B�����ziۄt.)� ���K���  ��t��tI# 
,JI)!�" ]"ݱ4�����y���qTv������ra
R���z}�/Tӑe��N�#�[o�ֿ||����١���?��z�zWd1b�Ջ�@�wK�t=�Ë���%ڃ�i�f	d����UN;���׼���.¬.V|>
v�;���~�>~�6-^��۪�0�,��޷���T��E4��}־<���6l�,��M�d�\�����W΂��29ml�[�g7fO�v��
*�N麭e2O}���_\��:��Ѻ�a��
=��7 ����`�|i�Q̶�+��`����ۻbf����{�~����"�{� ���K�$�.B����jXw4�:YY��)�tͲ��z3�Uj,��m��qz�%"�֗��x�V9&��"�To2� ;���d�YB"��PV���ɠU�h�=�F�lim���0])\�u�� �gZz�J�X����������n��^
���g�?kZץvͬ������
՛��<~F��^_�g�͟��[~�n��lQ�%u�������,��N��VE����w��˽������??�5�z�X�BK���w`�ef�g[���G���S�O�T��n]�F��h���ZMa����8���b�*=���r )��Qs��ec}ƾ�O�0���J�����2��)�`7�obg�W�Λܞ�~�I�O ����gn��r�x�ԡgg��CZ��*�o1˸|�+�V�XN8s�歘��7�S�E7H>Ov8Ϡ8�qHJ���5���Cv�8J=.��b˔1�fE�H��v�k/w��>,���Ŧ�8Q���0�F��Z�:��t=n�^7^��o.,F1�g ��y~�m���Bj.'g�|��>�+wR%8R��Ij0I�1�_np ��2��{4@����+
�	ؿ5�F�����[?�Ia�"��{TS4��fi���ٌ�ź@�j�ﲖ�݃󲻔t�U��NuIW�����C��$�/6F=c<��H0L��9+�1Ҫ�M��e�*��Z��.�d��O�RV�|�'|~�)�S����X�+���	�A�@�7t�h�g�G�團�����d� �t��^�nx3_�׽ay���е6����̴�����n�@���������,܅��,�r��%��� �a�6e7������s�#����Q�������=��7�hhU-�/z0���1����t*�y��7"�?rdU�
6%lʰ�I��㺎���]�e<p�¬T塾�����<ݮ
l�3?����yt��B���{�zoͮ�s��b�HDW�A�t��"�G˼���^^�hZR���5���/!����R���&��tF�v� ��d�%��?��u�T��R�s�g���WA#����~1P� K�h�����SB�xt���s)p#��"\���[�ܺ_u8F+ȁ����W���������vy����Xp4���lQR�����g�}/2�^9k�b�7�5���y� ��TR���~�oט���E�V��%���О���S߯�����o��o(.��P�:��L~�ӣ}���{Ճ`~v�_�S�O��\׮��Y�屼�qxa�q!���Q��ηッ�S�'�����ϐ7����{��)ݼ����)��*/��}A 5�###yi"���O�444�w�il10�K�J�G�G.�tl�I޿%$iH�A��$a�w�I�gB�M�e�9Z+T�X�ⅱ
Sf�x���~�=j��.s�U�����t�������㷪㈴��{�t�!��R�t�So/�O�Tp$w']N�|�G�1����W#���$C����ŀ����ME�WS����G�|�Y�[�<��}������FG�vww[��+���:G�z�A�°�T���=�����,��`�q)�u���U�t&����ۇ�(ޒ? ����&����4��#2*Wm��j
�WW�pt���)ьx�w^��W�&��o>��*��W��7�1�#�AlY��_0����&'��+J�[[O;:X�M���e�,֘[��n��se�Q	b(�
G����Ì�V��U��ߊk�g�A=�[Ε�1���ѺS4���p�0���K<N�������;��ۿ�ONm���\�jE���O�X2޸�B��@y�hz[|������f-G�^\\�����>���䖐��*Mnmi�655�'"�9��)����h��U���$$"�����{�X���M܄��N�J���l6�}	������y㱆�m��7^޵�M.z=W�^���^]�ϋ�[�%F�B��&��ţ���YG�2Ҋ�R>���;���J/��e�~\6���.�?'�-ύ��8��f��~b*��)vt��9�+Y��6�@��B�9��c���KH0455���I3G�LK�LJ�00�j��R���aT44�-�0M�����\�������Jh+*_��_�3V� ��e�S޺X{ځ��] �[#ܜ
��� ��q��*d!$(<��{v����G����v>4$&�㠎�݈�ř6b�K��y�R�e��Ku"G�'�4/[�m�e[���x7+�)���������?⇇݉5*RD"O��B
�	��d��o<��CYW�?�������F�Y�BfV�tth���g77�H�^�����o��E�B
;�m�����ĞO4�4�n�گ��nѧs���X��>VbR~Zy�'�w�A��%�46]1��W��JKgk��i�XX����|��qyz�:��Bj;���{��b��&��R�#-�aq���w}�=K۫?�W���-��q�C�-C8cdFG���(�^��������Y����*VNN���öJ������Ӏ����tq{�fw�;a\b�`���1#Af��8K�����ȯwX�[���8I��c*XM���R�g�1��ѝ�P�c��
fI#Vm����Y��-�F>B�k/E��ju`�c2�7���7�Kte������Ӈ��6�8�ﱮ3I5��H=�&���@tgq�3J	�������F}V��h|^�")ɨk���z���g�acoo�g�ںI���g�d�$Ȩ��Y��VV�)��k�C�&�AR�6�������:Z�->��SG/&�dD'�
�������X}�`e$A5"�oh�y�~�|�Bi��e�K��9+��uLp�e^��ܗ�/�H&�xܵy1��MS�Kn5������/Ok:Q�2�Cvv~�]
*��|(t�����H�_�k̎e����C."m�0Jw�33@M"v'��X�s�#�nh׾�#+\X���l�l��}��r�3}�N�:���sN����܍/���sh�fvUE�k@{(�
�y{e#q��9(Y�7~`��e�ⓐȃ>���1royt|��KGDD�&'��a��w�?�1��u��vT@CC��3x^J�G�(�єOC�_O�M�����^O�9��P�"��(Φ,��7�>m1�&�T�2�H�-1���R�K����D�z��z�;�����ֿ�^��#q3�S�,nC��(:���Ë�`��B.���F�o���Q*y+�0���~%U��)))HX'��1�2Vlc�j�}X ������x%{��ܢttg��ӄ�W�]�.a:
�C�<.)���ǳ9���o��}�~\�;���{���U�)�or�O±��z'���Z-A�Ji֛ݨ�-)`V_>�L�qy�ĥB11��$�����E�q�`��a��QE�	������xx�u|����꺀9�����}��o�V$��a���u5����e=O`���	�^�oa�V��+�HY��,��p��%=�p��O2^�ޠԂ`Fs�ʸ �|d��2�bϟ�H��-q��e��*�?[u��ݡ��KSR1��"��� �?w�8Q��`q
N��0�d��9j���C�{��DFFF`��T����]w�u��n��rYI����wж�� �&��f
9���~-U�������Mj����D����̙MF��}2F��1���z)��ܻ'3Kn�t`<'����f�]�@�Ysu�DH�}3�b2����O��/_�̸��{^ߐ�0��:�Dx;	��ݕtOI]}�����Ų���/�{C�V����m
����}���i�-b�q�^5~ZnS��Û0�:���ӝZY�&K VԒ�����@��b�w��S.�6�~��ш>UW��x� }�@X.�H����u���t�S�H��b��z�7��ha41";:�����"	k��<:� h	�oj4��"&F���`��0}ą,9n>MZ�/�=�ߺ%���,�	� ڣ��V���O���&�1�(~s����)��m?���R���X߸{�g?���������ނv�H\�>� }A�D���iP��6�Yמ�uX"��[muz�pE86�F����
(?���`b�BLxq~�28��o���:ܼ.�)$���۰���n�ET|O��mŻ.jh��y3,�[o�V��N�J��x.��X��a�x$���y����a��ک��F8�,3 8��zkvnQ���SjbJm!�+=CB	����|�ԇ����@qc�t�+Q3hf���V��Xؓ�����!ܴ%��y��r�������Ջ��sݶ ��&U_��"����������t��q��%�k��d'N㞱7e)�Y&���_t����t���X�7�LN*>����� u� �U�~��$K(<S�c��[�@ x� (�nU��&4�&L��4q��5{[g�����G�SI�1<�Jʸ��T8<<<W;=7W9�~Ǵ=����ݿ��N�06Q�E>���&��ѝ�`�=� _p4j�I�7���瘘��Ƒ�q�M��B�&��¶ߏ�V��;h�~K9�W�,�Ķ��N��BhȿdL�tk��$�X�%������P.[���B�>u?�o{�/*u�0��R�+���+~�jOA,��	�5�0������򚱩�Q��
������0%m�߷�V��)u(7E�S�W� 	��$�rq#�f6�cꋯ-R��mG?�Wz� >9O[���6q�A�s;R_q��CѠU��2��Kė-�-�G�m���R����6�,��0m���z���*�j>��nl �,�@�:�����D���deeĆHqR�2�Eީ�gbbHcgYXBfv���\{�~��3��1�ʧ$V��H���9j���!�+|������v��G'������bᐄ��|U��u��Qc|ͅ��>�(M��=<?�C�tG��!���_QۛI��ԏ�L�k����Z7����Rl��*XAz�r*))�.�|���2�3��.ls
s�N4������6g�f�c}�P\��F���G�1�o�����/��<�|!)���3��� r����佤�G�8|�!9��'��$&j��qdqN��rX8<V+�Bʀ��q�#	���v!���H��&���϶��LO�C�U�Ԙ�4�wu7�����Y��	��S����]�/l��ߖ%�$���-�.�Z���ub�W6��9�; ����d���p��uG4�z�Y��T�8�]���hۘ�����I���xxnx�_�Z�5.�o̎��5��J?�(4b�Y�4�Og�����=�"��_�g�G��}k�bYNNNץ�E��_����r��f���±uR%J4�h�<L3*
j(
E���M<�k3�����>�{�	-Y!؝wz���f�M�����j�%^�<��j���I�oe���o�K�vxԶ��(�,K@C�ihhڳ[��n�e	��'��#��m��qP��/�@?�JA��u^P�(����<_�KWRSKP;.�!�#�潎%Nod�;J���a�%s[Cπ����Ų��<���l��P��A�oA�hR1>.��>�{a���9�Ϙ�7Ȥ�OE�0�2��蠩�#HyZ�).Ge�f���W���<Ze���c�L�~9��x����nj߰�G J���TY�?��ͷ�?�EX��c��0�q��*-���"����kC����/�:��D�B�7Q�u� �"L��ʦ�R�<����:�k��躒ٙ�'Km���?����g͇q�a-�F���?}^C����9K����ab�'o���Ĺ1 �k84�̩MnW�Y�-d����f��֔ɨ޻�����f����+}�-�d�?~D�4kV�}W�7�,��9��j���S�0N7X�t�+��;9�5L�<8���$A���u�����ҙ�SF�t�A�x�����:u%��-��&wȡE�$T3�H���-T��6�as&�=��� �[�[�>n��,ȣ'�nm���X�p}�k���Z�b���ТSv�bK� �5��S{�|`�P�e<�^d����w�0A�/
$�m`г�����#Ҹ��4ג��`"&H�|���g&��YZ����JTn�g̫�i��X��2i���(졜ު	�i�ml/A� N<b�x�p�I+c�bB6F�UB�,9`������E��M�m||�VXؘAscCc� �]`���9� #��ѧ�����6+uڊ'��|���W^������%g�]41�q�q䡲�}$�H��:i�9�yG}`��2T�=z�So��?�}��qJ�6�L	�*kJ�p�[y�&Z�q
�d�UZ��r�J��(	���hR����$�ޞG7!'葏T�W4�Lm����E�U�g&�pX�V\��X��� ��Zi��3H*bQ������8b�v��0^��;�je0Pj�Eo{�kc�N�q�4>�I�K�y�>?y𦝰��笿�V��N2����<gc3������]Bs]Y2�(�MD�~DƧg�+#E�Hx�A�;�g��uXn7�st���.�� wqJ��]����R�1Ӳ1ǌ/:p��߶Q��n����v��B�"��y�j��x<�ʥ<�{�t|*	�5�g-֡T��{�g7����yF��C������_N��ҐZ���7r��&�Q��Z�t����z���	�d>|X��5I(V��bI�$q��~B��y��\^���Bb��z�n(��)̇ZF����}�I���>	�'��hC~�lA�i���Dw�1���WUŖ:����Z�4���h�M)�w�J93�2�!O\�'u�]Ƶ�{5z;�#��2=� �w���8SipS�]$��p8���ӧ����0"[�Z��s@�X�Qܩ��gv�~t�Q����1%����a]:��V�hZ���H�W��gv,�*�"&�F(tH&�)��ҼܝH�6k�$H���1��%ht���^b'�ثX �6#���=���ܷZɺ�2U�����z�pe&i1��S�Ŭ��"Urb�v�ٙi
�Ew��9�A� .�ؤ�P��܋��1r��Dh�N$�|�H��:
���=������� �j�/��Ic{00l'<��0���D�8�q��ﮬ�v�:��I�I�ɻZ�Ab\Lˊi���i�G�p���<)�oę?�Ԛ-�Lt��J����AM,D��}�j�"84����~k,���p�|3,�Ml�"|@����}"2��� /��IH����je�=�;�' X�l�V��3�Sr��H^���=H4�m����S�8�,mx�~ t
.b��g^��	Z��s�hth�¬�p�c��B��������4�v�ʮ��<��gl8�?�a��}O�|��j��K�MAx-���@�Ϟeְ6
�E}���6�\���]Dһ��N��|�#K��u�?�H3��?��G�<B��e���R����*N�B�b)�E���I9�x[jH�,������'E9�Gl��1|"�q�zI��o���F�&�ȟ<͏�ؿ���۫�� >4f}�� ����ײA�M��/f��~�Ԣ+)��?z(��K��ZZsb��C�C��諓��]M����|.^���.�e�s�x�~�/��� I����F�"��?�*%ǉf �Qi�+s�`EΜ�w2ӂ{>���9�Ւ�&��C
��-�Q9��*_����]`_�{!s�5����ك�0|4U���T���N�5�Z��ftaf���V�K�p �@�ĉ�U#�)�ںM�`���r�{2#�Աhnf�=�K$70�������A�ժiu�Z>G��W��'�������F�%+���������J�eJ��{�0��yH��(7^ML�W�ePh�'7H�q63��pM*l\b�/����V����/f������*�� ��t�u�����Me����8�ړ�\v]�^�-�zc�͇A9�,�D�����9y<'@��V��7ExPO �}�~���4���Z����	p��Eq'������7����S�[KAg�,5���^3�gn+��_<X�Y��#z�0$a�p�a�����e^XX���@ �^��i�T�g>�"i_mA�����ģ�~fc���/���JZp�j`�������Ц��=R�.g��ۻ�!�ܸ���-��,32����E���� �=2�<D�!T(&CI��4�[�1	fsC��yv���û���[~�f	�5i��DQ�ښ�;a=|7o^;?=\&y��̻�Ăd<uGGi�l+%�ĳ IXFi�4B���x�RW
�u7�����}fD�7�Y�F������	�棔R�W��׭4���e�)>&�<���aG9G y�`Q�ƖQ�H;���B�"��ZQۓç�,OR�־�SB.Hy�8Y��t�U�#�[��a���NO�|��}�/WW�����o�������'2uFdAM�3��S{�/i��&&'q.��Tlmo�����n\M��J�Zu��;�B6�u�^��;H
Du��s�S⑽�$@MU5�ZrF�(	���l�<��� ����}e�/��T���m�F�x��e���3�h��칬��xhFT�e`u�Q�Rx������3�m4==j���7[�	l�G� ò5��8oϔJ+[��|�����<�2> �]]���D)�!ss�SE�2�E߾�;���V8:9i��%����><T41a!ƽ��/4�������sR;���Nm�N���߁�a�;����$�c�����Z���~��=0܄ǡ���rN*����U1}Ђ�� ��Bj�i:<��HR�O�M#��ъ9F�ddF��`3���V����{59ƧD��=�����7uw���#�b������53|�T�ם~]y�/�6�K�2.u���=�E�����9���|�Eޤ��B �zd�G���4}d��x����]��#'**�O��G�T��� ����yO�X�5ɯ_��K��u��`�J�OD`��iFF΀A��.��6�o:,]ԝ�F�ZT_qCV_��:�U=f�ɞo=�;̈́zf�)T���k�+��Q��4�Խ����&���w���I��}y83�_)G0/��Me��q��8��uͭ��`����Z�*�������X�7i�鮿~#3=�j��J���8�F�<�yڪ�LG����%��<3_��H;5���F��h
����h6g�:&�����`�ZZA�^&��$)8�Q���'�k2d���}Efn.~��F���Ν���Pf��7�����c�q�Yɻ��]���O��A9�0V���+~"m�=��JeS�2䃔���ʵ��7�4�	T��F�)9P�����`! %CN�`����8$�����9��u?A�������5����1�tD:��8.���k����Ɨ��۾�����y=�)�f��:TЈ]��}��
�`�,�N��~���N��cL�y��|[ɫ]�4I�ݥ���'��dc�/�g����k8ҹ�s?�yؼ�0��d,�XG���c��3�M��o��[�{DU��Ə�Y���/�]�h6�8rD=k��#%l�7x�D�}��Hm�gӸh��KUrR��eԡ��v��'�p���'1k[I��b�ج���:�20tI���ol͈"ox6\]B�0H+)5ŕ���
D����bXSn�{~�3_<>�j�ɡ��\U�,D$}q�������1CGǻ����u��] X1N�-+h>@�c�
�j�����Ī�St�l&?~:�z�=c⚌Å�m����y��Y%Ay�+_&��6~-c�b�����ϣ�����WX\���u�t�b�����pٟPy�.`	
����m���+{����s�`k(~Lh��Y&I�fJ��x (G�1�"�=���ذ�am�����c��S@�u�ٚ*�r���{}�Fw?e��/���?%fz%�q�{RÍ}�q\]]�n���ѕ�@��>KQ�yɉrJ��������yW9[+��ë�i�4zfp˭�����Y`�e�2��3��`��y�p�Hd@�AG�N���*�p¨!	~��.�J�wee�0��}ʗ�e��pzG���S(�bb`��@Ӗ�A)�76\�2VN����������y�z���Б8����ŕ���&C�L�t�-����\]����0�j+��4�}莵�u��N��T1ʵ�"�'O�#נ�+�kkk�	�-׻^��e��Q�8�?��U�j��:4��<Cy�lI?�ƻ��ƛa*A,"�-1ǚ$k~��~d߯FZ%Nu������K\�]��ԟ"��oq�o�!#���f����NK�E�3]��~"�E����b^:_��#F�z#.����y�~��wa����[a��U!!��J�K-zl���oݠ�/�:����f�P^U5�8����t�&��[�_�#��`��"Eĺj'd1n�d!C�̶|��c����3�Vx_��m�����"�M�PJ���k�y�*��!�;���`#�?�c	��O��~���ǀ�*�,-�̥s6g;x��ރ�����h�wa�g�Dx�����2��ҙ� �ŋ�$�1����Q ���R�U���++H������U�����K�)�����,B��s�+K�M"�H�j$4Is��j"�lk�)�@�dh�iz�w�2����I�|�ꥤ�ڗ:ҝ�����c��c`����(E	h�<��~�g�r>@g��rT�A5�'�y��^���~�L�I����<�%�\�ϗ0���R�57���
�`;ZP����c�1%�O*1�/Fy��A�@
ZpLKK[̉A*����zP���"��?vK�����[����G�h�;��H��+�-�����$o�8�����*$K�5�DC'Pa1�Ç�7P��%�	_{��&�r�g�ܷ0��/HV��!��:�~I�������r�������g�~��!a����5?����.�q�2ջ>�¨�V��D�����m�~����y�:�T�n�ޓ�U�Pנ	���G)��5S?g~AA����[O�][\\K� ���@Ǵ?C���/�Ǌ2"�q�oߚX�"����^��d>Jta�;�/#m�(�K��i� �Sw"������"`�O�����嚹�4��Z�_z#5���T�ZA��FW�l��U��������Ar�|�8���ct��~��e��gk�)��:�n���dA9� ��
?W�GG�sO�ٜs++E

�����mMAx;��ӳ۳-�Hm���S�����z��ŵ��;��W3:����9@��c����xk��r��������Ѹv�žZ�N�8Imsh�w��V�槃!��Χ�Ls{�(( ��7J�_m~t�������w:(��� �#7u%񀢢�
��V�=��S�g�'u�����8���r'���˨��-���]�Ȩ.K����g\��;����A�Q�V�;���ώw��~�B��������VQȤ�)��;b������.Y��㧇� �O_2�ޏ��ZlfHV.J�OŒ���~3��ƚ,�$���Q�#JXo���
��۴���/9���4i�,�Lf@���b닔���	��l�6��l�|�4E�k�EFF>4���.��o�ݼ,P����AZ@"u�r�7��VR=�ӀN��c31�쳮���%���y� Ɔ��VVQ)1i�Z���w�1���R��N���s�� zZf���x뫾��+L�K���\��c^�7�&��aL�4
�$ο,W��]m���x�Xx��-�B��x�@�uǯ���7��]����_{d��Ccy�W�U>�:��72�ԯ�B��!^�TO���j���9��8��@gd=&!�y���t!p��~W���q�З.�"j���W8���+}��S[a��_��.v&��x�^�k��=As	

*-�>I�_c�5>�9Y�P&����{������4,4U5���)6&��A6>Z�$�|��X��e$R�u$�;�m*�2��	ȟO����o��3M)����v���2�y��.��0<��K��L R8[7�s�w=�P�ZZB�&�� x��Z�ȺZ�Z���zx^��>�zw�ek��q��+�䘔�|��w|���85'�PR���W��������5�?X%ٜ���y�����*��>�"��٫���XuY��Ae�"*fd��6��\k9O6b�?m���!rW��#Ğŕ��o��_�R��ն�UR4j�g��{(�����88��b����>S��9��G��׽�Fڻ��|���߶�e����� �2U�ϵ9��[W	a��JD	������h�Pn^ޫ����Qs�yyy����!��!5���H-T��폽*���_|��������MWW1���!
��<�ƣq�Ν�g�`�Z��1M%�Ji�${���T|r��j��9��Id�땃�C�&�a��Tk�􁴴�2 �}�.�it�n~�����J�C�@��	T�����8h�l��I[֩�ڧ &	E�7�����	� �NGۦЁ
	�߁�rg"��dM�C�Y�|bb	ΕC��Ɓ��:�z3���L~w2�࢞���GЅ<�00ں�ad�-xު����z�B����<�]3
����=nh{����w�5��������$~�4�����[k�#"���M�Dt�ӡ"� ���Z��*m��_C��8����-���+�g��+4��1i��rt��K7�q3=��X����m_av~����{ݭك�I�S���8��;���Mk��f���m��by��^�������~����Q�'��i�4���h3T�Ԕ+�[\U�gY�7=�M�lo��������4i[ND���`��z�Ff:�:����K��8�3I5�W�}�Kt��~�^�{�OZ�
s5ş���U�$Q|�`��(�~�ao����n������4r��&|>�n���7�QhXS�o�}�!88��N7(�}V�^Ó���|��
lh��.!A�= 6�迗���]�{��Z�)sL7�$��\�62������������Y�U�S����Y��+-S֩	�i����A�g|S�/�z��ê�\��w#��1���m�H�u$&:���E&��S��뿄��Ctq�-�ۄqW�Κʴ�[S��)_��'#@�-��Dy�W�[	`�<��Y���:j��������?��(�DXu4t>M�ʿz�:Q5�����Y>��� `��0Z�����0�Q� ��(�����-0�	�X(G��H̪�Q^iGL$$���Pk��B^��:؎�Pc�y|XY�$i�~?|��}��K&��ۢ�v����=������hk�C���tb/wX��v��E�K8E�=|vvFNْ3Bd8�\�
<�(0l'ܨ�}����`H�]�;KʧN1�&��.
!��<T�y�{��P� �h��|?4�j�����h����#�U�l'�ǉ��$v�f><1����P��.,X_�Z�����"�]��jq��/�:�0|)/�i1}���6��'�c�M�@	3$W#%�,�[�|�WN%�M[���K_�	��W>v�ѿ�ee�'�da*՝i��v�gD0�����*9}b�����K͒	��nsh��lG�:wux4@/�;_#A��B�V/\�]�h�~�{��v��t�u�|�5GK��/��g#bG�������Oi��XP�D��}���lh*6��y��׽:G�J+�ʥ����P�|X�~�9�X�����fm���#I_��*��m���999A����s��R��P/��+�.eTN�W�+ڧ�;�ƺo�L�#E.�t��{AR�,�þ蟄.ܵۺ;��"�D����Z���V���JK�J�a����`���C��β#���a�.�;5��&���{����@�Q��s�ďꌽ#V dpo���ԩ ���x��Wc��"h���}�I�|��������n�3������A�����Uϟ���<�ĜB�������_��Ӽ�,&v�%�UZ���)��*so>3�$���U�eP�`�`o���9E`������F�ۖ������G`����p��" ��|�~=��_��
�DBo�PY"�,f��0�N��tCq޴�$�e�gD-�����?����q��J����?dV#�X�9��ߠ{�(�����ⓑ%�X��Ru��I4�m�8_e~���Xp�Ǖ-�(�{��(�	�|�tg,(}�'�jH��p���z��O�S@���z|c���1KH�%ũ���aa�J�y�2���}�b�(�Sf��H��������� ��n��TˋM���W��Yc����|���ry��S��Q���_�@[�3�]�>�b͈_]��qT�
y�ܯ6�z�h.��V�.��=<R���U�B2��o߾��=DMM�W����S�$4Ĩ�|Sf32w�dǀyh�ó��G�LrΜ1X���2�Y��Y��~
��<@-��oZ �SqeuwCȰyߥA4��EfƷ��)-��7��IE�Dr����r��p�S;7�ӥޣ�=Օ~�k�u��������C��HO̭FJ�ۃ?�!#�q�<��0��v�	B��!F���Z,��.ǥ�F�q��XL[.�pjȽ��3��Wc��u��.���g�� ���hllm|{٩MQ����?o%�֭8gy�����-h�U�ͽr� ���c8pz�S�����KK˙ GkS��wj�h�-�1�笡Q�ѥ	�w��Z9�����!*H�L�_7l� �|Q����q��%���'WR�`�-����=ci�4j��V&&j��N�f�ȡ�V�*��Ӽ��y��4����m}k?�k����fH�
�r��͂#�7�kCy�H�F�������t2eeez��U�"s>V�"�����(�)*�@�Q���[F�i��fB��B��Ӻ�J\;W�eת���GV�j�>8m*��~#K�A���>C4��J��SA��]v��g�<&T`����@4�����H�x+J52�ii����o\	wh����N�κ�'�a�S\�R�uOu
Q[�E���U�U�:�n�a�2��|�8�:��?�t��D����Ƣ2����,*���Ɔ�Є�̘\�v��VX�H��d��m�`����^���e^z�Ե�p�j/H��ǪY�m`j{9���jYY��G�W"��޿���-Z��5f� �0��Td��; ��;�Ξv|��&I/��b���㣳�����T���Y��=�qߤ紁*	Jf	��8Τ��儘{ҷ`���l��>o(�o`do�>5��j�M�{��K<AH��������2�ӧ8�>�*hR]��a�������	��Z�������.113+����1�eI333�
�����C\��ݟ�	)((��1`��A���j����q���
�T�<��Pd�mߞ4�+�6�x���г�ӗ��7/N-��Ð��P9߯�f������5�㇞H��OP�����5�b�c<��]Jr0.=�E��mYt��,W����)+7^�� �#oz�@th�
A���Xo�(�2�N|�U�  ��$x�懡Эɰk]I�1Rנ�����(�d]_�����;�5X�14�[\� ��S@��pK�յ�����B�0I�U8���`�u����~{{�?#��yb���KШ����ݹ���*�����T��ڍ�e��)�N���hmm���Ȉ�!sۚ"����z�$t��2�}W_}�� =��_o�"V��ĺ�]X}��%kB�Eæi)x���f
Yq�H�g�h�ּw'�*�V:�����W|����߭��:���(�U�:c��ܴ�l%�@��O%�7�H��l�s�Tc�/��Yg��g�Z���炌L�] Ș(a�%8�4���<[�� �H����n/ǘ~9������������ܜ��X����ˇ-��7B�df�'r+����L2�e�����_Ŝ� �"!������~�@-��>�1���ɐ�����������uMgaiI��{r���5�w@�0�C��uS������?~<3?���3tk�0�����+Jʘ��R0������Xu�BO������TV�S��	�f��P����5}?�m
��QuUֶ�р		;�	�O�=��:�[D��+�탶��<���|�Ǵl���Ry =�C���^��3m�:G��$��@Y���Rk
�6&|Ym�4�j����P.#��i��jO�����K\$�N17z+��;)����T�ޅ��Z~�K���ᣔ:l##�=%�y���@N�Q��/��|O��y�6�(^�,n��APX߽{��ty�N�eY�s�ã���Ƥ{f��Ʉd1�C�F�`��1|��XO�>��ݵ,�!e��R�w����<pHOvO��l��]��[�@>$v���������-L�u��կ������f�M�/O�R��0� �T�@LD^vDS��K�a�m�od�F�t����4?Zz$�m�U�8�0����G�U�ׯjy�s�L�j1�k֍�o��G���q#4Oʖ'����G�E�=��p�2H���-?���Z�L�~�ז>���̳";(\��O���"��L�^hi��0�xˑ���
&�I�% ��*��T�/��Ķؤ$�ɨ�����iy���-��A���3���?~�7n� �>�1H�LH����K��_Dn���2��k��TpUTnе6��}�M6OS@SYsJ�_;��|�E�^{>���͆�����E*5N^�t �wwX��p�3hS�Q��9 �/��n?6�҅Ylv��N�5�G�uW>Ҋ���B+��[�����|�9I�);�r�-bq�5w�T���_{�Q�����;�&έU5�����x{@�f�Οvly�T��S��ĻE몕!�b�j#�D ��'f��TLL�����(��2Z�TQVT? Q�['�[�^_�	����s^P
~�:�����*����-@�,��:��I�RC��c�+��캶AJ�.	i�.鮡T@D�)Ii%�a��R��;���A���?7O|�����d-\é}���u�s�3D.)�t�ʷ����5;�(I���OF��z��%�������<��s��b�HƙR��W�o��1���9��'��8���P�F�&&���`7�M���h��Y��j��F����衖︍&�/���ǥ�����y�x�-g�Ҋ�ޓ�FF?������0~��0:���D'�]����@w�uLs�!��z4P�Z�tm����5ϧ@�����;C����?s���
�3[ZZ*�T�����=2ؖ��Ҋ@���*�-MT���ݣ�������-M���d�r�p��|�%>�^�u:]>�t�FKs�,zW���	7�h�l,B��;�8�9'���PC���1�3o�,C����󽎀fT�c�ЩO7��Չ�a�΂���i��!�|ɰSu����9��v�o��q9��U?�Ed�D����cX�ϳ��X��#���ȯ2|j�{�VI`���f�z���R�F��"<h�>���lEz�g��ذRRR�F$�wO�q?�l�~)-���Qu\�:��P��3^�����m�����4����ZO?@�݅o(%�Ջ3��\"h��H��~�괫p�����ZM�X}%��/��\x� &-w��S��){rM�W�1����������Z������sx^�D����u�v�?!�v�!�W����p �w4�cA���~���h9ٝ8��ԃ�����q�[�i*m�͆�����:�xӫ�7�u�����G}Q�{��c��O����Ĉ�Ӄ⃂���w��Ξ6p+��+m��՛B���O���z�J\�6M�G
4��X���kn���"S�&1�9H����?عI�ft�0���Ɔ#`5��dJ��r�����Z)	����3/���������44H�h߰j���Q�|�7޳�Ҽ.���k�n��������ۭm�3"��v���_�a�/r�ѷ����<b�H.h�N�2��DUͷ9�B����@87�I:a���d�b�>2�}:q8s�Ւg�_[���RI3{� �f�sI2OzĦϺ��	3[-qw6=I�T�`@@SU�#��NdoH���G��9�n���{̝�0Xc>9�T�4xcqpn��||�܆�zv����	=��[Њ,��;�� ..���
^��TQE�7((�J[q�?��!������o�IF����Q��mYߠ[�����'2�������OJMݵ��{��5m�{���|<i���t�9��_������i�H��$;{$9aюl%��v>����"��}�	O����f�g�߮q�X�k۶��ck�'O��w{$�2ǭ$��}[G����ڥin&���x\�~��I�t��9�`<��כ9����#Tt剴�l>�,j��9=����Iӯ���1��sf�M֫�4�6��{:�o�5���9·�rs�����o��zE��AA�(��]v��3/��sto}������x9֛�@8VN{�l�R���6}�3����a7Q�����WOܵ�ʺiT8��l�v���ʟ	��̓���8ը�Q�_��J"�INƕ��!.�G����]�+�y��o�}����b�(-g�������g#m?�dv��AfG�je�a��������c�Vt:��ʮ�CݘN1��5s�n}��2{�|���;�眮h����ͦ�� ,�Dߘ���ҍ��o�گ��dVX�ڛ�.�ѷ��d�@[����v�Z�nfaR������4�S�99evc�}��l��-��rrOܯ�ű��H�??jeeu�A'��4P0]�̕	�T5i�kWv���&��Yt�ft�0N���w|���&��
�P7��T���yO�u�F@<$���������4�K�C��6m t����)���{��'��ħ�qBc��빯��G���f�4&+�.JL�PZ�ܽw����=+���A�uoѮuӁ����i^nN�����B���0s�-�ev�(\��X���t􉾁l��T���9��a��7�]S��׷�2��FϽ�v�Z����\��C�B�	����uY��=��k��/�^��J�Q#ф��g�^�L�4��]0U�۱�Ap���)�]��*�����*O����n(k�:�E/G�K�1�v�ew�!�����u�-��˙��
�����8����dH�GW0���|F�χ�����QU���f�;e?�b�9����"��z89�^�kt���\�y'�Ī��aa��Z�pۨ���ZxD0���& M���?���8�Ag�;ts��rqc^�8}�v�����?3O3f�]~CM�IЄ̈��/�=�8��{l�!0Y��EJ�x��r��	=4�73=i��G����B��;��Ѵe����C�}<����޻��t?l��PSu"��n����V1$�S)k���=���G���{����hs�>�0�χ��2{�o��w2���6a�|5��Ľ�(��{�SqH��H� �%����U��~ɔg����:>9)��x�BRw7>���x��X�VʃxvL**����Qk+����`ʽݞ���~j�s<�Y��]\i��dOiA9��[�c�b��fsy��׭���fL�%�C�]mY�q�m��Q��k;�-(>�����ɈSɨ�5��n��(��ʶ,Z��ڽQ\���/�	[���߲pcj� �(�h�?B��)(�����20#41W�E�K���B��py,��6.���P�t�H�=v|�M�sM�P���T�D8c���1�7�Ǝ<�T�Rr��`�Y\�	$��q ��	���}�Ŕ���y��Sĉ�w�8=�%��[��gL{�o��'�����&��!����̇.|���8�c������H�����4�{�\]]��yQ��J�z����--O�?�5= :�sq;�^ҳ������?2]�Ԍ�C�UV�����J:u҃�ڦ}�6��� ��+W�U���m^���y.�=��=����H*��6p,R��Y �У��Iߴ\��Jj%���v��/П�&GZl�U _�|���S�c�C�ӕ����O7����q�tE�1��
*a�O��c��<؈X"�+ҳ*��J���I�ɴn���m���Ht����(��'�N��Y*�0�5������>�C���B8N�E���@�~[�§ ��RPP@��l����	bV�ٲ�9�=���"�1��^�L0��q
�F��^b��:�(j,&�ԛD���R�A��l9��퍤{�F������`yY/���Ni��(nMU�Y:��5L
���w8��(5_�j~w�q���h��p�6D�8�a+�&q;cH���)�3�� ���Ha+�����K��Ԏ�P4?Vг\	��Rw����%k=gs^Tkb��ϥ��^� x�Qf�Ǳ���FæWB�������q:��V��i0��qԬ�F��)(���\!0-"&����J�����:	�Xw���y���}�c%_�� ����M����)ǰ�eN9]׎L��+�V�~F�0��,���W��~G�|[��ɗ�r��G��1N07x'\r�:��1���-q�YCS ������.B�ӷS ��B�ÞEsݢݮ,UV[V$�L5���F­�(�5��R�.A_ `�9S�v9v�WZ��,*G�} �28�zh�L�����}7���4�x�c���5뼽��b���W(����
q@���� �(�T3ߺ8t�����O�doZ �C%���HA�#�B�vVx���ٍ�F�=��RI|F��wnJYM�<�.ծ�N 3�䓲0���miad�>��b^���^��g��<R�'�z�¡I�}!�'���B񎾿L���?��D�.Ui�yٖ���w�Q�|����aVZM�C�k��3����6?@`}�c�ӯ��4�3Jx�:�|����߭�%��j�K������lp��G��޳Ñ�ΰ��X:<��&"P�E��6�`�x��̚�֥ͪ��p�pޫ����;�sʟ?����E��nZ��&"9)���s�V:ך��gR�V� ����SD�u����2و�(3�IǳJ��u3+;�x�S��ϟ,���Kr@����z�_�Ƃ32A~FhѾ�qT��ф���w�Tю�������:N����"s����}�.#�.G�X�SI��hA�$�3���-� ԃ�k���r٠o��cA�-�9����tv�LY�,�Zv-�}��4to�b�ܐ�����Y+��e-߀A�̩D8�����O�ωOQ5Ǖe���%��!���U�E!w~�1 �u:0��%���`A�wO��Y>��u��O�OW>(�(K5�/�/z�N��!Be�|�t��h,���:3�}��f뇎�5�8^G
f{{6n��� �-,�b�� ���g����Z��/^��D� �K��Ug��T���j���CL�H��c��m�~��T��;�S�5M �x�K�E��[�3GWI�����3�oi�]k�����(��K�)��}�+�}Uo��ܽ)0IX�Ǡ�q|w&{/֋���G����c�ښ=��&V�0�)��m��0tά��ߣo�>�A$(A�T$
�Cы����x��M4������$���]�:^��̈́)=�*Bf���2�	���� hv�?�2X(����)�|��_Wz�=����cI	5R��
��0@�w���]a��<���=�<H�a��s��zo�۲м���+��NL? ���n^��]�	�Bk�� ��c�~���gG�H��F-K��p��Zم:����N<q�/@sNŜ,��Zf��z>���?��KY��ڷc�}�6=}�$�F&�d+��V1���,����U5a��I�����B�/5�0�*2��������uc�U�{�[e�^Ă�}5�e�|�L��FN_��2&XlF�t��u������>���*�}�'@�Gٲ	+�9Y�]%nȓ2(�>���؈|n��pp��Ѹٱy\�̌���x�D.
!l=��mk��]��Gj䢲���L�('/y�����y;��	Q\*6��M���t[ �O�t�z3$C��H�d�p���_!��ll�6��I1V-$"���s���0��e׋r���%��0�z�ذ�G��-x(@	�W�αJ^��O���n
lF��n`�<.�E $�^���-l�]���y6��[}d2ez�j2}�\�\�s�
Ec���;����W�4%��_����b��&���G?�k45'�j^��D�����g���V���R���ϗ!u��/���.a�,�WM8��.�	[�0	^��R�>je��z��T���I���bqq1���|����:)�%h�.����xz����ެ�P�:R#����]]��Xd8l����i[X��jZ����FRYl ����H���qh��s�4�ʡxb��xba���u�;J��Ⱦ�m��G�_!�"]qc�KN��E��{#1���#E�o(�.�n��3����yY����%�R�)"fV��۟S|��>��Қk�^<�R����υ܌\=��X�K���$��(���ˌ]�F���|j��Sb?��ݎ�أl=��Μ�o��5ۑ�fEJ�9������ܲ&��4 �� ��llHAȃ���Ζ7K|���nei	x�cKKv��%���8�{j�]���Ҍ`�i����I$�?��t1�V���>���T�6_��ݜ�����۳�k.��0� ��ƭ�	���Q�������|�z�[�cE.��Є}5U{��N���)�!�~}:�����nq\R]#�����e��S)������a����-1���p�y�
a�R�r���;,��|U3l r�9���*�O�Ý�~ݛnb�Iz���z���e/�sz��%�-���j6,�w�u���!ֆ��fE���"��A���`:����',��!�εX��*y���7}�<vE��S���8L@5�Ʃ�9�����%˞p�4�,;z�y�8�v��t��
�����H��֦����x"�Ŀ�Z��%/�����ss:��l�v��_ۚ��a��d�����e*DƸUJ�W7���.������[�����P���˫nپ����ܳZl I�~��-�ϲ���~�Y9��3Hs���	��'i�����;4�ӻ�2�ڄ<z��{bZTpii�u�&�b�\� ����kՀ2�S%�����E3��%�А �NAA���Mߊu�#���%w�0k@�>���p���Iq!f^į4�ù����]~�xu��ub�@|��k�E�W�hÿ�Fv�җ]8�uZ��?���4s(�.0�-X$��Vo�}�H�^Z-턘�����o�?e���;ψ�B�+2L%�6��{��|~�ӶMX ��S�6w��5I2+����L���5O��S�g���gt��9����>��r�Q���c�ҙz��?�X\���v/-N�Vʞ[K'q�,�R/|Q[}�[ɧ	UJ���Z~����66>���>�H����噰�A���u�����z*$u<g/�a����9U��ڶ�[��3��4�Kj��!�r$�e�� �de�I�3�~.�;ZCCVK��`ʖ`�4:`7��~^��Ҁ:�W��Խ����){�JR���S�������0�K�z�ėr
�+�p���Rp�8ѿ�ym���&���O�7�I��^�h�V�������&��}��?<��:<����8�Ժ=�����gwJ� ���[�^Vx�,�������?-	�,ŇZK���}�Qh:(Dc/���n��8"��5�;��5N0".�U�#?TWSyyy�l)BGu�A�S6���ԋj���-����/J>��W�PMP�w��4���
w����!�7!a��EL<;���]��O�G���M��D�-��dFOci�p#�7�t~'>-�3��iW����c�'��H�R���t���M�a��W┐�I� *���VU�q)l恚�V���/�:�N��y�S{R���}&��#90�E%����Ԉ_޵7e�.%&)ġ�R1����t\+�^&Y��Q����M����6�m��)e����CK�4�I:�~p5�Pt���w�æz��)���%����*�ҧ��d���1�k��u�c�{p�ڌ�H��&�׀�����*T��d�T��ƥRrI9)�а��S���a+'�P�C=��*�w���m��3��
ӡa~�.��}�H-H������������nSw��k��3,z�B�7��k�Vq��:�t�H4;m,��0���MJ����uy��O�q�H�����1kuX��x�70okt�,�ǧ���ʖ���ͥ<pVR?��~{��pw�(L����ăɲZ˝2޷��w'���T��9R�?*D-�ϰ��c����]"|g�A̭��I��Q�/�	d�A�:���ul.���\/�)y5v8;4�����_�\���;1d�C�m&�I٣��Q�F[�+����."�<����?�a�d�U���I塜ݱ�N�oR�s�O&]��%�E��j��k�(F3�M���mL?�O�^ܑm�u��:�b׌�}���k��R�%J <����KŴ5�,�Χ��HǞ���U�Ũk�򻛻��\����9پW`�E\�)�1�uNk-3~x���|�����	���0��}g`�-τfM�[��&�լ�F�-/���	���/��DE�o��WKlw�t����TU�E;>��a�NսC��Č����^a]�,�es[���:������5{�!۬�}��L4� �(���́��#;���ΌJ��'�B�ڭ��d�|�( >![�o���!��5M��ׅL�
3� P/z�bnA
$���I�p	wn	W��y��@9V�K�-�d��k�B'.55�QMkJ-ʙJ�L�uf�(�k5�A����)���ӭ�t���Ũ��h2d�'H���1�T
�^���)��3~(J@�22��`�h���������,��k��I6׽ﳙ;�%���z<�r��F��{r��P�#��7+m�>��$�|R6�܄D<k���bvO��e�Tt��2l{Ε_H����v?"�H������bg:ɣF����(wW<��]6����ZJ2^7�TzmZcbp���K�c^�y��1G�m�Wt�^�]�yߐx�J���/���h�����)��� �my�b���?c弡,i
.�@�����"�G�#I�e�:�y���A���r��!�����O�7$�#��H�L��������Ԑ�9���+�@TM�/��Ě
Gd��k�Vr,�w�%��V�Z���G�RH46kΖ�E>�=�V�i��+]���Ӂ�ܲp��_#_�M"$���*��T	+F,y��p�veoi��#BnY�h?.��!�K�g��i��QUs�SQs-�����l��T~�W�Q�|���u�,=���0}$A�m�52i{��5W�C3p2ᾢ{36_鏘����{~�L�;r#�DC�U+ӷS�K^ߐ��\��x2�����l}��+���G܇��"J��l�b��e�������<�|1��<�E��T�r�+/YM�Ƒ�
�kF�]��0@Μq�8u��K��Gܞs��E��S�	������5m��*ߓ z�����J~uv�7MD�7<�*�* �!RZh[�z}�$�}J{�N�G�����JĞ;ȏ�!��R�~� BQ�����=F���{D��]�:������L�i��鼛�Tq1[��#ED�L�;?{����^���v���<��onKS�FʥG̾UujO7z��Ҕ�l�v��x�'��=��io*:;�X�X ��w�%�)5_͗�������u�$\�-��[4�"�h�A�\8�r�����whep��ܷ@�T�������}1EM
�V;"�#_?)��K�������*�(��'D����r�#���u$�W�ݬ���xS{)����mv��w8L������H��cg�YGN���qG]g��	
H�uA���@>&$��N��
��uJ$e?c���p ȮO��+x�̈́ٸ���a�o�I��uӐQ<�j(���]����FGk��utJø߹I���J��!B��6���թq��(Uu?=>��y�Åm��)Q�jq�Io�ב���o'�#*r� ��3�W���qun���&�6�G�A"5�9?vҩ>�:��v�	Ju�yd2�����3h�юV�C9��t'��[��ʦ/������9MXˉ����=Bn��د�}�c��7hP(�e0`���#�� rs<�|@==:u~9��#[:$/u}�T���h��>)�H;���+&�Z�S5>\���u`��'�։������sxz<"z0�tJZ�fm7+���"��9,�̾��O���/�"�"� ��V���Yg����Y��]<-B	��I�w[m�����4�6eY�~����A�w���ԍۀ��=�v��p�����B�v���
��a�A�CE�P���V_9S��EB��E:�!�,���s�4�E�>] U��tD�2S`Aq�(@�W Ջ�P�|��%�|(�]�OW(_ݐ��+�z}����Ӻ	�8�v�����_���b�W�>���;F}����'I�:�?�VR~smO����>� 0���Ǔ�MI4�5��s�H�����q�0�]�J>+���~y�|��k��/���'Q�V|���R���߻���c�(#����A���j�ܐ`H�[�������鱌2�%Qΐ0v�|ޅ���	}�w�I:Dt̕�S�LǾw�%$
��E�e\g{@����ɦ�G�In�q3d�z�)�e�H��4���p�-֜�g�=�Ҍ��#,Ι}ݺԡp-��L	7"���ܱ�1��f�z��$�y�T���٥+�}O��aa��Ӆ��`H� �C�z<���ʅ�u���N�]�~WMf�l6�Y��[G��-�����Ƶ.�!��������di��^Ak�m��~�hf��:Yr6C������a�����_��c�a�@���C�B���2���F`_���{�~�4[�Lf:a0���Z(��d��fωMɸb�Y$A_9\Ti�4<��D7rN���MqIq9x6��z�9<��^�+�j>�:�R}H�^qb�(+�ݾ��O$����bO�s��^H ���tW�)�z���4�p� �?�:	����Bc�38?>^�Cpw+���j�þG�v��pH�qڨ�R��Q�3���n��8v�0���>�����_�ޅ��AVI�I�v3��W�:�A8��hWZ�z@�{�
̮��J�8��F�Z� 4��UywZ(b$�ާ��=�st�<��}m/\��o��xv�������>���#8�n�K�T�kY|tㇵ)�z�%-���;��W�畞�O~�#C�(o����Xl�Lc���;*@���_D�ʕ890���f%�� ��	��ٗ�ެW.Y�gƂ�������5�5ȯ�x�#����@���������y�׸8�A���6>y"�M���s�`j.��}U�<3db�0��T������$&y�/a����;y��E֓���r�K�Jf��aX���x���aJ��J1=���lc�l�Ӄ�s��+����άC��t�V�)��6��^������R�w�G�G5$��-��%�<{��L(ɚ:�1+٨��7Jn/�ۏ_�EO��Em�ʢ�6���>��9��(��pg���j~;���Q=�_|n���6�&�N��@P1�È���0v�lcT�Co zAL+GH��@{�X�B9�	�߾�vT�HV^��8�+y_	:T�e�b?����iP�Р\]LJ\�8���w��*E���w$ɗ2��&hMԔ�M����`���`Z	��j���տ%�.$Q�qW���̺��i���~�4ZˌK��m��W����B7�R��������<?<��X��֮Y,��z���DTl�2�|B�Q�h�P=�H�w|����7`� =�ܾ"HO���S���2|��~��ҷ�I�w@s��T�nNn��"����|wV'ȶxZPc�|����IpJ�B��0��~����Z����`׀h��7aJ�E���ޖ%�"_��!ucQ��d��L���pr��
`���Ԩ�0-.���%j-h��i��ʺ��k���WFo�L�LW5O�M҉m�/�3�T(��a�>��h�ف�Ehe��,a(0��z�携o�z��K���#�eP����o��S@PB�ʎ��)\%�>�		�(e��	�gKu�S�Tݧ��5x��(����7w�gYr�k7��`�$�-6��j4%7��M�ě��G�r�0���h�_�\��($$��*ʮ:��giǥP�L�S��=j����;ymk$�78�⟜�8	'���Et����<����zR���M�`�Ě��NŚ�D�z0��Q-�e���_#{���Ʋ����G޿�M Z�ޭ~ 5U��Xl$i�h��(v�ss)t�l4�N$����Ƀz�Y���3>��,j�n"�{��9ݝ'?�<PV�I�3��j5t�˔�����3��TLj3��;���T��b��������a4ߥ*�ޱW��fP�k��%��q�2x��?&%����
���u� t� k���\�Zx�iil�
rۈСh-@Y�>��B�O	����!A�����y�<$j�:���p��zV �}93��vH|�����$��_�t�[�� Uo��g�-O��T�ri {!���A^���9�D��C1�s�a�`'��*٠;�ldW��0M����,�}��Ǵ��+�p+y��O�,ioW�����fx@�I�}bt3���V����8l�W�eϠ�O��>n�Bt�@E�S?�fj��y�ة�+}Ι2��"�!4�囙��b�S���j�t�qj�y�I'QY�v�⮸�%S,��;P#X`���w|� F�tG��'��6w�륻�j�&R���ɚ Dp��
]�r�+Ԛ�p7;��̫�ꟕ�Dj�P���Ϧ��z|drd��A���=�O�p`���s��D}�^�=Qx<��A5_=R7t��qm|gI�s����d�$_S��B�S*%��B��>�k��g��~F�Հ�~&����`�H̋����v;�̴:��5��,"� @��pD�0� V��_X�#E��)8�h3�#�pW�P�2�X�^�p_ma���~b@�-�I��F�bA$���ֻ��/����7A?]ې��|���Qq@C��q��Z]������go�o�mV��䀹U+��9����q.��.$ CC&y����-pC�JU:��M�x��F��\��D �'+����!�s�K�6�l���l^n��2�<���^�_�I��d2D!�`��z{�&�z.ʊ������!��ˇ���]�c0�f3�s^*�N�B�qE����h�̊���	JǋtO����h��NeE�t��T������"IY��2�P"B�[�Ow��r�v��2�"�����??q���s?.1��M+yiڬ����uEz<Ж͐_�w\\ м�	622��ی�<��=~���hS�-&��V�H�T�ID|3�k���gO+^M�p�w� �tn2(M�7�H�c�9�A��1���Plb��b�q�!��w��j$�~o8~PXK1����C���my�`T�&Wြ�'kM2`h���Հ,��� ��\8�IT������X�z��u�H�[nK����I9�s����x�R�\��wX�㎱�]V̩�g�r�B�	����PK�#�^��YE+S�w)����JNtfTߨ0������i���a"zӆ~�9��QǝQ��� �7}��A��2%J(�c

b�N\�6��0@����6�����L�XlC�؁X�z)(*_:
Ln(u�v� y�.�r�l�I�
���_��� ��5�B�k�	������/��"IW��аTj8���B0u��&�Թ���^l����^v:��A��)�f�L:^���;�	�7�F,VO�x�*�u�ޕ/x?~���[��8���3tB)a�e:m>N��m,�$� ���&�q��U�� ��fv{�]2����lQ�KA�����^	�^��������F��<�G����\�z���WI��n�U+u:�ª,^:��ן�x�~�DI���� �3'�ȕbh����1��uV�ꫨ*2�.	X��K���tw��sZ
,
�X���W�y���H�Ǣ���&��"��n���x2�.�����M��a�����Ah��{Q&>�#���=a���q���Avᾄa��*����H��A�ֻ~�B���N1{.�	��"r�
D���vd4���N������v7���,��<�PmO\д.gI�]0�$c}C ����ɋy��yw)�H.nn�j�'��A���s.�tC�"]:k�r{���ӽ��F�	��֥���F+o�¬ÂE����9��� My���@Ǭ�3��\Yd/T���� �..#��u����}t��)&pP�x��[�[X	й���E�q�l@qaaK٩i�q)j�q�����irG1R��b}����Q�6R2)��+�
ʩ�/^�p��_����Ύ�����`�y9t�C��
Y�+@M�����v�J�vk2B� ��(K��/9�IX4�F��)��{�봈{�DH���P���8��)�}���"e�=������1�ӄ�"�/]����>d��{�E�{�-���!���7u��sm���c���]祐�Wq&pc"ҾD���Mͷ���UY�)E���0+�����p�&''g��a����GcC$e��%�x�����>c��Rc��@7<7��m�C����8)�E��R)F��^�M�i�֏(���4;M�U� s�%�8�`�;�F�D�a�ʵ�k�?�}�A���4��Z�p/B*��_D�J{��D��kӏ�䧛sm:+`p��1���e���
Ea=�4ȫo���V�W�Q� �2���ep����Lz�lt����P�U
�Cq���Jh�����ާS�m=������!�6j��Ar� �"3m�&��L�v�b.��Ez���Tu�:�����׹a�ʈ�:��(��I47��a�yi��ì��Q�Z|�G���Y
���kW�|�F�*�P�h�go{{��ox���i[�HD7n�W2��D)�b�
��rt� �G�M�Pa��[��wN�Bg�83����#WQ\����,�LM3є�����M��c�v�����|��6b �6�X�X[=�*g8z��Ά7����� �1���X""i[a�����4�J5��W�g����x@��+��f��aD:�}H��]={%j�J�$������;��2���ip��Hп�`M���}�x��Q��蟧��+͖�J�	��me@ ��:�.ht���	�9�	�.�.�Q��/�7�^uӚ�պ-�.����G�o�Z�Z���3&'i%�c�\��`J�&J�q�W6U��ɪ%����Թ���p���!m�� {��m�4&3��`:RQ�ǱV94l��m�r t�D�ldѸ�S��Su��i���?i�_�ZF[�׷�Ps3��}�
g&D�M��^��|z�f$���?QBW-��$y�~��%v_&���R÷*�`)[^!��{v��'�:!ۂ/0�0h�I��7'����M��ֲà8�������Z�xK�GvH��s�K\���.$g``P�ԤB
�$$P׍Zݽ{ȗ�1�NM�_��k�D��dv�x�����Fw���><T@r�w��
&P��霻CSR��d-��1��"yq���
D�kᎤ0~ݬ|%Lnh��7���dCk�3}�pj���z�����y��
)��8C�����&Į���E��~�yF��Õ`_������8ǫ���U������@��ih@�����;����}:.M�i}}=G���z>%:�q����ɱ������w��	{'���sg�9�=T���i=Q",H�Ю.����֖�piHa��!�����d�(-�+P�����I�xN�gW�F8/��X�zR��k�|Q##�+�A��"�J`#��_���#�׃D&�������[h<	�4˔7	>���������QB+;�v+.W2�F��Ϡ."""h���� �[.ήe�&%Q��<��PQ����w�.�]�}''��㿞h>7y�k4V����"��?����^)���G	-4Ao��䏲�^�WR�bna�b}E.����Q��R���~��)>)�Y>��c;� ���xw�#'".qy���y`Cؘlgo�:�����V4��A,��ob(�7#�À�\~���y�ɠ!Z|���)h[i=�����Y���W��?�|O���6�zc�p*��f��9���R�����o~�A�^����]�X\B�VRR�̰f�R�xH"�ul���S����V�y���M)�K���`��X�������H!��]��.��w�F���̀���޼�⎋OJA8=m:,&"t�&9쿟p�Hh�p��
��8���$0�h�5��#"X4��	�EEAC+�׿���'
�8S�%Z��8�`�Ä�����ݫБ��$Ѥ���˩������e�Z������~h�͗4qm�����3^�3{�V.���f��^��%�I��َ�t#>�Y|l��Ի�t���׭瓼�'��<K��L���Oњtx~덂��:!�/�������V^o�4K66c�d��~���-n�o����r�~�M'%%���߅�b��XF�1Ա��߅w�ͼ>Y��EWY߇QQQ�L�x�|�:n�����D[!����7�=��#B�`v]V���o��	T\׊k{�\�O�xpٚo����A�[���<8)�{�l�h�lG�w����P$��/c.���ZeM�mc�1��V|��ߒ�W<��d<���G3��F\��t��N6{lb�7��4����~��M>��LZ	�JO�_�-���^�͗��:>��k�0��If��%z8���I�?���@;�����4)�[TQq{�q��F���.MП?���_D2�J�s=��Ƥ�oa�{uXX#33'���G��TӪ�S��ϟ��\덧_�َ���7N\�Q322����Q�6���?�qC+�.��<[̀o��v��1��[���%ݞM�L��f�[#�����R���,r?�p|x��P�8�������n�	�7������K�����-�|E�=�up������6�6�|֍���M�s5EC�tG�>�LMa�Sp� X�pdl�����xO�z��'��˶���\��[|�x*�׹]���@���^��q�[9[Cc#�gNa��H�F��R�h\�H�l���դ.n������R{��]5ϧ��?�����4��@@Um��׸N4[<D�c��?��iV`��2Dz�4Sn�d�����~�0��ZȻ~�3�/)��=n�˶�'e!���9`;�ޕ,da�>Y-d�9�*?RLl�g����\�{w�|�
#��_ZЦ7�)&W-�,�������Ao�ͻ#�s@J���{���. ��UZk�����a�}���]�9��fg}��]a�o��9Q�� e?=^OO����@̣B=�L����v����2�)����%��+�q�Q��&\5��P&�|j����'[m.`�˾�M�f�'�֧j�2dR�	���$P����D[[P��7�ige0�U+	A��ׯ]�4=�3���lqi����������sv�嶶ʯs�q��D��}�c4�')Y����[HuCCC��,|q�)������릑��me7�����ǩK��ܙ�ii��=�)��s�� ����
�
K���@�WǻU+��@�A�|��>if�;N�<�����T~��^ȋ�y�I�Зe�W���⫝&�����Ew�Hƿ1�љA?�ߵ�s�y~�9�/�g�Ew8U������Vw&�n�v�l6����ߑr�$(}v����������[��n�x��� ���:U���nH���K���ե�y\��Sj-��l�t4�t��'��,����)��I�~/��������fY�M)���AFV�vz�=�&��N|G�`�o���=��l�>eȰz�����P�S3�3���s�O �T� Jɝ]M���&�X��X��<1���bO��_���z��M���c�+O���9�ק���T��ku�H�_i��\��bhh��qqn.[ƫ���M���c�v���|��j�'��F3�`�OMѯ�G�����W����V L[[{Rw>�� �s�~%��Zt��߿�?@<V�� ��E���;ou��w�nmBB�B��dm!e/���%ٳ���N��Qdٍe�2f��Ԍ}c���>S�u����9�9�y��9��\��z�_������md��h��:� �E��^ա����/.�!�!���3�A�ف8�p�:i����lomZ6ň�	X�������7-���)��$.�:v��9z���@���Md�|��dd2�趻AY$ '���#`Q�����H�HHL$Lg���(��7\���;UH@�_bs�) ��J�Y�o�~��D���K'e��9\����
�Z�������;�w-.�����/���^�k��u�Vb��C�%|���b���Ì�k�AN���JOp�l��t�Z y1�j6�
B5xR���a��F���&�-�NBB�A0%4<<�$S���"y������������Hf]U{{����J��׭{w9���R9�� ��!��5r�s�����)�q����\�
.�r())�V:uq1�Ʃz��+ܛ���i��'�՟���Bv��-�ZZ^���|v�]�����������?��Q�-�_� "����$��=`�IcQ���nH�ڞX�$O��`�Dr���@���+�Ỳ�mu�Z��� ݮ�i��AL�cQ���4�u��rJ��q�5(�߁9�
���xLmD�{uO�ٴ&�������o��Ehá9���eȌ�)m80$*i�ML&��(��;6��
���H/|ОZ?�j����$��!��<	(x�o4�{�'@�O=ĥ�V�{�p!��{����8�U�����J��e{��K�������@��K� ak�H�&j~/����o������n6�rO8U���J\�ʥ�H7K�* '����]	]XX�"ձZ��|]�[d�/_�<Uq��ѱ$�;;�?�MO0%���1,�HX@��+v���T�E� $����AX����NK�Z$+������C1���*$1GIZj?�`�-�7���IK��/_ު�r�JQV���w�[F��\�G�P�m����q���	��!���⎄�s������@�睙��&q4�����ÿ�{̨������ $f
}7׼j9F�@
�_�Mt��ý���'2��%���- �d��8ށ�Ds<3$smk�hjj�W��Vd^���J����Ar���,d )�6�D�,�^ɱx��� ���� 6���.P^,��������lI��lu������PB��~�H��k�pK?�W~G]kZa��xKH(̗�B�]�,��^@�7�~z�����ђ�Һ���u""�A���Z������7�^ѳ�2 ���Q$^�-��4^����柡�vn��K�}�	P�G�u���]����?�?Q��� �����?�i����=�:������Zɋ��T��M��}�}�ξ�u����+��8� Jκ���I�.�N���ځ����c�bΌu3�SJ�_���d!+a��������8��Ͱ��?6���'���mn^^X�m�ۿW��~�b"+��(��|�ĵ��z�۫r~T�?�"ۥݰ+ՠ�S��S��^	0�����X��xS'�"��r��߻��\H�Ǌv��w������7��5�>f�7�	�LX�OW���3���Ԝ/FWis}ȹ���B'{���<��ia�F���Aq.����s�Zp�v3v��d�p�^"����k�y�L�ut��I���V�(}�c?��IG�U�Km�;�ַ��_J�~� ��ȱG8�i�r]x43+�oS>++�G�7O�n�BD�]����#��M/Po��F]�<��`�P7i��!vk�1"+�޳q�dϫC<H،8f^ű��e�����M�Փ�z�,��4YX�U9'�]�6v8��Ү�r��ҜL�N�;�J;�_yyЭW+���%=����J8]�t�c^��x��>��_D�?ےrIǧV�3�r��@WS~M�&�D�V��F^��@���%o�G�f�p�(�6��o��>J��:�ٺ�mR��K���G�^���=:��#rS]u�B�fQW�O}l.�f6F�ȫ�*�{����]2��V�:W#s����9�H�.�1<IH�<����#����W����,V_��=2��[{�������nt��N���ȭ���t��C7r(Q� ]�Շ%&S"�h��K���2�%��P���M�	1Y���/��#l'bq#�<��eE&���c�V^no��*�190�aD�辰�o��	V�;�ؑ�)���!���|��1ޞ!9e�G��X�v�hIA�U�B�j�׃���]�q��Ѝ�8�2^���� Ka�ۡ�B��֑�ٙb����Ɓ��m��V��+�/P�f�,E�ڇS�){ߺ�%��#�g�t;A�0���~t&Qv#�\�2CQy+�6iv�����@{����|� �z���j��^{�3��88�)����a��iᤗ��*+�y���9ƶ��3Tu�Orw%��{��#��t�}�{�R%H�Nl�%\�Ԫɭ��Y�c���3rxY�X�ꊼ=
�G��$�����8a�HхK� c�;y#�11t�u�����#��pmS��D�{~^����G�m�������Ǆ0�!�Fn�d�-�m}|V�;��	�`~׽�#��{#Y�Դo�������>F��U���)���&񗌔KMw��f�����fFҝ:���C} �CyLS�6C+�&�.�Ӽ�).�1􆄵����KC�ڊ����n����]X�2 ;�K%V���8��U��O����T��`{��U�f~�V�zd�(|����s[n�A���RH��b�������o��Y��#�-�JA�"+�TVF����5vy�b�r�,F~��GW!W�J��cs8�bp�sM��7M��
&L���-�~ߴ����!-��ɢ|ٜ��'a|]l/��n^Ш��
>`�.g{x����
e0g�����LR��4�	^��&;��@Y'yw���������K�?�����!��]����t ��^��H�:hJ=���o����=v��7/��<���ЅF'c9?brqje��(��0s�ied�&6�{Oɍh�����HԾ��Z7i������9�,��OO��P�I\2��Q�m��B/7I�U��/�f���t�)n�P�'D2���ߖF>`жjY��Ab��!ޒ�hlҐ��wU�7r�����Ϭ萕�[��ަ�9"Q����I�7�Lc���������)��R�f��M����2Y+H��Ss,Q��,���
@��υVB���4s�<*-b�U�6��&�)�qlާ(힏!u٠s"�����vxh��Μ)kG7�1A�����T��,<��I��K��W?��a� �X���O�u�ǃ`=���^锔�p^E�둝i�δ��;�
.�q2�P ��=��7k�4���_���L��%%�婝O��W�\�i�|��U���hIY��<-���ڊ�����ɱ
ۅ)L���8F�'%h�����8[���\d�Cu�$l�
���/��0Y���i����D'(���?��ھye[���H��In�a.����$E���K��(Q�hk�4�5~,B��653b�^����XO�!frTVvDNp=@s��5��Mcg�+�������A.mP�N��s��Ϯ`��Л�|H$`����VS3E���ńJ���ۅ^N+�|�2�T��
Ё�!�}JJ��'w�6~�. vFxnp6AĲ����9KokV��q��T�S�c)޽(C��ut�+�tA��ܻv�P��ϱ�$0�2��xM���pz�VĨ����T)x!�X���,��; ���䢽}��#c󓼨��i
��0����D�%7�����,3�
��S%D�Oq~{v�.��.u�J��^{���R�ڹ�.������sAYHy�k�-:c"��}K��gU.�ɜ��p�0\��wmR�+�B��l���2�>�Z�.bP�}��9؆-L���T��qjn�J�]D^� ���%qfnlhHU�
� ;zI��`m�IW�qO����fk�.��J��r�τ�W9�YL�N 	��8�\���.7B��W��Fq�B�|5_W�^cr���q��ٱ�Y_�c�Y�:W�vt� �z'1N���ஃ6 ��m�(�!��(�\������+�k4Ϣ����5T+-��!�cTr�Ā
*Y,V7�A6�S,r��iJ�-S}C}+���
L;m;�GU��MVV�l�,m����%��&�I80j\�Y�Vx�(��G�@8#�_��">��d��Z]��v����Z>*#Y��Q7����%��$�e��/�'��{9�wj;Is�n�=�7�����U,�(���(~t�T�� $Q)�>Y<"�s��^$@���>lXN�Fe�iX�_��-&09������Ҵ�ŸCN/Ç>�5 >�� �V��zu�dS[Rxİ�h�+|R{m�x.H�d��B������<�=:*����ZkjY7xP�T`��Xl������c�Y�nV~q	C0���)��^��t��*%͒e1|<�T���an�}D���cB�� �mu�jb~C����xx��P�sp� ��G�����RW�[��{��ʄ�F	��X�vP�Fs�-��ѤT�|f����C��d7��U�V-�}��I��\!k�>��Q�0ny�.��O/��<5��抣�QE�ؼP��n�c�68��;�N�R�us�G���_�r��|{� p�Ip�a&tg�+�3��Y���a󾺯�s٪xU+��o����P$���u-� ��v�0bF�:g���s�[��PCFta�E~��1^�hA�1���ګ�qG��K<r�`*�g[��?�f7b)���r)��3yke<�M{Фf(`nmA.i�#w����Q�o��,�#(�hN]�\�2;� ;2�j*�U�aoXX�����D`�B9&�u�{��x���Ģ��>N�~^�xE�m/�k��g�4�'��v&�	��@�����~1��_�J�z��YbJ(���A#۔e\8Ne+�T�[l�\E�]���Pt�2�f+�_�Q�Y$�/10_��=хھU�b�|en��h��k�Ӗ1Uq3��W���k(���+���2zT�Z^����Q�i�6ꔯ~��wֳ]��A�4n��A]�������/��:���կ�@�^�~�)S�V�����L/���|���뇋���j0���|��_�:�(�@�_`{�3�I�y(+�k*�ZP�>�>X��<�b�'���|+l�nz�ƶ�q� ,UdC1������	ߜ�w66�\�x�/9!�Y�)�׍��̛*ᛄ��9�>��v��9 70��%��#����	xr,�YP䙔_��U� �k�d]RU,C�γ?�=��$�hK������?y&�L!K� \fcU���x}b�!R�m~f:B���F���z�o�_��G�%�F@��Td�C\�[$s�`���עy���6n1A�'���}���^�蹅��)��=�Y�C�f�����P�i1S�w���,�$�F���� ��L%�����
&G�3��=��N���D��.�S���O6OR�yx�x��󘸒��$w���9^ƿ�q<�&�i��KR��.n]��yq#�m�O=�����]}h0�veW,H<{��\C�sr����7�יV}��b��HYy9,�0)���,'ehG�X���Yh���520`!�9u�@���]98��-������O?�6
�(CL5����M�֋Pa��J��}'l�;DwY����yߟ}�zNډ����ɖ�׳�[گ�5z|�9y��/1t���딚� `�_+y��)2�om1�RF$}���U�9��#lw��Y�DIc,��>������Ѣ��6H�[2b{;E��H��nA�'�{F�)o_fį�q�������$�T��!F=��N����ff���ώ��Џ�by .�A.��I5�cƃF��t���CX��]�'/�}c"�"{B���}�	i�������ɚ��؄�MXX[�����LH#ksu�oL���P�8ÁߧO1�6Ap�M�\9OP7��ce���v�/��nn��]�lO�=l������Ht�Y�u��Ɵ�\�<hмͭ )H����3�L����@����V7�Я��I~�����P�2z���l�������$X[����g�B$�ǟ��ZS�؏���L�X�7�n�y̫2U�L�>��\W�:�fSI`6?�i#�r��Sh�3KI��mH���ͤź��诧�f4�w:��ف�r����m�0������P����q�(O����y#Ȼ����y����?��8��:2؃�Jy�=ol�EV3#�SNThgA/3��?[\���T�TLKAp�B~��)�`�NtEd���Yߔ>��!�"��fWn�(����.���Ȋ�ѺԹ��GG�d���r-��~��k�㝔�C��u;�%1��K1���x��V"��^����G�'�v�828����iD��IB\��M/���޵G�.�,"��tn�X7�.�x�b�P��I�Ŏ�ed~�D�Vg�j��J�G��,�)8���kʲV7��4���m�},6��1��0%>R�!�����eꂕ��Z��#5�K������Ԧ
��j�n��'3��":��	�9����L� sZ��x2�]a�׃e��R�w�����[�i��=Vv����o�"����1u����7�L��KŒ1}�]��eO7gZ7�����]�W>C����-Ӯӭ��ھچ>�/��ˉ�)�mR�HFF!�Vb�~ա����g�9r,/F&���s���ĉ�m�W�W�D�ȡ���
s�R|7���U�����ӋȟT����'Cf�4~eM��=�ƞ��?����u�R��1ۜ��6��Qg-�5шC�Q�C���a��5����gc[s�O��`�R��Ӯ]	3ӬC8I�ф�\B��9��q�+ʜ17G z���QE�2D���_]yM��T�JXA�!�geXw긚�Ewj%��|��6eI����������̧���o�� B���|i�y��v��w��XӼJu�8��i|��8�k�bc�>���WC�O�qR�'sTg��l�Hc�Ձ;��q�ۯ]7�a�}'���S<����5�M����}s0����Jz3r���ԗ�\7���N��� ����l�R4���gfԔu��Jg�����IA V|�	�[W�;�$qĚTK+��Q�/Dy���nBZ{�����w��Z+Ԇ�z��exS��m�J5,�{�zYB��5��1��eå��H����\F�K����a�K��O�ニL�<�O���{���ܼ�W>�3��E�_)��en���zW�GT�����t$=��>}*���6�S{Z+?Kp#�bw����xͷVL|�
jM�3T[�,�[%���|�k`��URjyF���ɫ��������n��@����P榺	�9VV�ܴ���c��xFB��+#�=4G^�\�~g�-�gv�A�����Q�&������WS&��'�-��'�l4=�AK���uok��ǫkc�ܚ3(]�zN)�u�����R>��}V����s�����&�0b_Io�����U�,28��J���[��1e����Ϫ��?�a�U�8��UEn@b�W��~c90�`$R��%�5��Ss�v�1�`���z������6��)j��6@���05:U��ij��Px/��{C"��ԛ@V�ƄJ�r�J�~��[)�jA'�k�b��Y���i����Ȼ�Қ�yZ>�܊L��٘�5��J�Y3�zi]J��!eED���M����
��k��X
W�6�
a+:f���߼d]J� l���؇��[�z��ՙ�5�?��3���?���[�^��l�m_"}�a�9Ⲍ�h3f��Z޵V��]���.@O_�����o��E��Ka������P��*���Z-�6��`ˬ���m!הI1-���,Z��-x9��n:���`S{��Wa���=�wz�o�w�Z�	�D\�&�	9�%jǓxg����c��O����&s��K��m�`�#I�,�/��=J�M���%�
�!��n�mu�:%z���E�{SJ��]�m<k$���Lz�����ٔ!��9��\r��.5��%��d�HBL��^�r׋��a���<5<�D��n�pv��������%p�$� �G��~.�N��~.�@e�g�8W��k��ɚ\t��?�)I���d���6��Z��]��4Abϯ����C_^�xw���+z��Hg0_=c�̇���u��SC ��z�P�06n�I��� �\��鿸�,��)ÊZ~=��RCR@����+5*�[_M�8����$E:{�A���P)�R`�{�+4�� Π����+V�X=-�o�<k;Ģ4�^��Z�L#�
��2���1W*v;������-^�Gf_ono������Z��.��^�4,T-��T'���!����SKoS�L]��뒛�.!��������wJ���)�zT��B����/��{F���w�Z��Z{�dW�ͺ}#�A��0&a����b�2�Ѓ�q�gJ����q�	('>#�YX����Kq�8�~������g����V4g�w�t��=�Ԝs��g婵K�wѠ6?���>3p%���NC��W�9���j��Rɇ=z�
o9��P~����A���/=��kP'(f������p4��Z+�fP�N-�L苼��峒�0�8=��H�����ȦSR�56���7�g�3�9x�X���48a��e��$�%�{o��j!���%�6�I�G��_5�~� "\:�O�i��*/�̗�v�w�~b���	�!�򦌀�f��a�$
-*�&N�85��&�i��]��k�R��;��_P��s�g��3Q�ꦾ���Z*Ka��S�Pcq�;��g��wecv���⚅ˍ^�׸�q��6_IL��b���e�ҡ�?ե�Ⱦ�׉�LHw�ٌ������_���Mv���߭�3��y�>Uf�|S��s��J��������4{h$�T�r�_��Z��{�Mv�h�a{�	�'5Kj�Բ�-�6	)�����ׂ��}�2��`Q����k��(���7�aF�k���2�o��z��7>���I� ��gm^$5%O�7d5ߞ���XpF{��Tx F]ߔ���2���wޝ���.A���ŏ������A�Z����}�Ҩ������I�G9پύ*X�'����=Eʍ�2*s(+�1�F꒙[��T��	J�EIZ�%ww�{�b9�s�P"mJ.n>ߕ0�M�A�rU�mO�(�����/����n/��5$�l?���8�q�������'������ ip;��_u��#��2��lGX&�a�ww�9�m$��~s�x�w�k ��ƒ4ʯ	AY�kBd���P"�pULz�|ؓ��į�������Đ6s��#-~e���Vs��eB�t^�U�?W&9����|�9�n�L������k"�=�~әZ�P1f*b��t|-��fX;%����i�J��{7���[.(����@��,W�4�kb%��t�0[�#�CM�����^ݑy�V}VljYGR7������ҫ\��2�$�z��gLԴ�'nH�V*
I�ʅ]��-�U�9i����ы:�2��r6g,��H*��e��"�dф QZ�����oJ�ۓ��z�B�"�#��ӷ2�ʰ�t{BgeWbWf.�x�«��ɑ�:k����l�^�R��M/ƃ�bJ��\F	)?��� ,�M��E|�*��/'�Ԉxnnv0�mpgOVļ絗��-�����^��R9����:�lQ໔�}�`��*q�w|�qG��sj��fblt5U�@��Y�߈�%u`�"��CÔh�_�% +��u�#�#_}���N��~U�
�`g9��X����Wt��2��p�0����v��G����ڧ�X{3�Q���FK��F6�bx`��⢖�8>>ْ�W��4L�\hs��a���c�tw�{u½���^�,�c�ƭ��#�a���#�!m�==>UT"��MB���Ms8'[�p����}	ótC嶧�=o�|�yMi��ߎa:��oU}8�#fO��VLac�GQ��lե���-_l���J�S�X-.�"�^�Z��������N�Ў�R�9�Y%�q��*���H�=q�A��A��9�n��z��m�-�ۉ��k��(S��у"WA)P����:�@��������_W�2p��;�le�+�����C�6uv�O*[	�و���,�w5x�o��}(FY-T��Q����-H����rV�L�$���.�[�k���N��C��Ȥ�l�m�>��ΡP��p��à,7P_����V���������q� 2L,�� ,|½��@����\���aΐ�$��AČ�8|[ڕ�$h�?6hޗ�^,˜�v徤�BmKn�!��|�Y�>)������:�X��nj֗�{;jZ�wE��U���|g��9���S�i�����t���e�1Ce���D�֊���z��I��v�D�ɛR��䫊E�r������
od��Hc]��I�$�O�^���Lx�{�ea���y��B��C�oӚ�9���=t�������#Fw��t�\tK��� ���Q������P�h:χ�,����P�;��R�ڑ4�ݩ����4�	o�A&��r����e��o����F��X�� �T<ol�>��M ����EK�<�쓊QJ1%�1
��r�3�}��.s9�<#����D�Ø��� +W������$�%P��'��w�^���pCޘ� �w+ ����`�9�qг�Η=)�=���y\	n�`[D�}AÜwa�����a@����	�J�>��y5-��s�sfZ����2/u��.S<t�[��h����`�����d_��ծ��ڈ����BF�.%2�
eAdY`Đ��>�(}��3����b��R�5��;w7��k-��uL�mk��$?h��h5ebM�>��O�T|o�Ƙ��+S���\=���d��#�7\&*˼��;�2��޶��S�q���θ4Yґ>�]&�w��s�T��<��z�|hG��tX��u�<Ay���������Vl5��<G�l�F�:�C��^H�8��w�V�0��O�/A����pUϳ(P�0����痤��
��˰B�&D�W���W�w����Ӵ�I�ɳ�o4�W,�ۦ$K�ֹ,�F*�m�*�a
o�&߀�>�/��4��"m3��峰oТ����޼�4�8鉽P�Fa�T���U�,ь]��?u�m��M�L}��X!-�]_�ˬR�����G�%E��{t���ց�ۣɅ��n�``e��MSp�MM\B�x��'rsfX2q��E�,��8�
S�f�y8��Ɲ�q������sؔ�Q�eI<:'_��Cw*0��v�`�l�y8�p���UK��r���:G
|����')<�L��ei�Dy4�X�(��.��"�#���a39HK�	%KH�f���H&�{?�^
��U��1�#-ށ��]E���|sP�H�wd�q�����/����.��y�� 4������]$�B�h����gQj�z�������D�W�*%[�w���{'�t�G2L-I/x��*��I�R�J^�F������~'�݆Q����FN�EH�,�C�`y�D�����:?��2� ��r
`5z��8j�qL]��{�t����/� V`��y���[�>��{�V��)�,�v	׷�l�(�Z��Jm��4��˽��[�nke��9��tc�t9Of_�}8T�N]|6�<��Ĉ������g�$�2 
���9�\�ݮ3���\��-:21�OV���O_B92,H�#��]~��������'�T�k�a��5r��s	��dy��O�sª�U�h2Dؤ9?��
�I�M~/���
d����uOcܻ��7��>~�&K��$��sצTP+M�d�ӺCO@ +&�?CYڙ[9^u�Z
�_eܒ/X{;���^�y����AP@l��~=���̳�N^-��'�,j/g�  �����Q&�A��&0ŗ�0s��Ҍ��!�!UҺ�k!�]J(P4�� �W��$�k��D��^���q�@�G�W(�u֩��� X�y���Z�Tb���I��Fh!1m!|���v����LZe�z��� ͑RI��S?hm7���huml�@/�UaF�I�������3Y!�7kM��0 }Lw�3��3�
(Yr���Z��\�l��f!m���V� 3��^����L���kX��
Ӯ�Zt�V,|ߊ�P�,.jU��iU-���sò�΢u�����7�<<�ME����@�8��@� ]��f"���
�����ʰ�I~V�ՏL�Ab��ͭe��l̋����YXҊ�$�{�zpT|�|Bg��E�3���$L=�Q׼�I_ma�Ν�E��v-�+�L��/,G�-�8�rD(�1�t��>�9S���i����5�Mȋ��Z��S�\����>㗄\YC�Y;c���YI������'= �G}���o���k�<�2�D��x xl���v�}:�(��-_��X�bql���̄mTJ�LJx�}la#�Xh9�	y�]��$7^&	�s�2�դ��y\MVc�\X��lH��)v��`���j��(�..˩9�js�I�bA�5ҐS�����ʞ���z��D����0�oL���(~�z3H������@"��u:�z�� ���)��L&���Ǟ8I;��m� ��B@%'w��+ep�W�4���ׄʍ>~/̦t�����P����u�u��y.x��wh|e��m|ᱧ�#��bR%�Lmq_�_�.�MM	�v��-�h�m��{F3`lh[��G�з��TT�ǈg�b��F����)�[�C��{c<V}�~�APS��Z�e�9����E�Kӽe�Ո��<��11�*_g���B������D�7�ʏp ����sqM�&g�� wJ=�ܴP���uj=o���S�jGw�g�ϻ[�����g z:Ee�p)��M%�Os�6�#;�-���§=��>�Vc&�l�=?�ޮ�p���4�����Юák���R͎�s��[���n��m!t�d���(���(Щ{��At��恀q�A��� A_�c������?N�U3��ZIq[Gi������5rv9���m�H�"eũ�q��c���`F��K����.�h�п~Hy�ҫEbL�ܩGM��Č�Q7^�����_ (3/<�O�����<�A���UB��1���q��g�����C7mKPP�K�y^�AЪF߬�����j9��R,t<��?^'��נ���V��[%��0�1�5(r ^I������-��yd��E�ۭy�G@��4j�5
d��.Ä���<��iσ�n��Kc��YF�AO�$�Z�����Xs_t��MB)�l�oZ�{q��hu俼Uλ�4�f��W�͉��_e�J��V�l���y4bj6�����1�S;�. )_Ӝ�?�[-�c�()Q �������?����������juA�y��~������^b3�!*�@P�y�g5���_�zϴ��u�� }ﲿb�w�󠬣��*2k�c�[�f#���~�4x-6��A��{2p<�@�^��E�zG��Sv���!�:��Z�\�����C�a�l�.����Ѣ���Y�`#��uVl�L�}�?�V�����i�A^�hs�b@e(�6�`j�Re)ܶ{riݣ���	:�b�h�՟@^�rs>��}v�T��]]�▬}���h-ڣ�����b �  j�%ѩ�ԡ�� J?a���IT<d��ۓZg>�gW�}��4.���/�:8���i�2�������������sc�^2������g��v�vt�����
u�mǌJ�۴<%z�p��vP�|U�/�t�p�HLm��~�Y�f9�;���k\;#T`�R�s��彘Բ&����Z��Hd`�KZ�`<����~s �hbg�4����86K�$,��&pK⣟ �-��_%D�Ѳ�*t�hj֫\���I�}#��p��pN�ը���^u�V0ף��S��u�7峒,��7r���3�-�֦v#�v�?\	�^�v<I��~*B���)�/K_��L���s=�sB�;��k���y��".���_��l�`�F$J/r��M��2�����TU�u��o۴�ɲ�ImV���ފ.'�(K��a]��d�|����:��X:��,��T��T�"��[�kd�ȍ���O������|�xm��o���`�i��'���O�4�^c���C�~�2띨�����?9�U��z,�s�Z#�9�
n�-h*�������q��,�@�8���Ԟ� �$n�A�(N�����/�r|"8ySp	U&�?�:&8;@]@CW1�ml��
"�xhxCLv����W6�n^&�䱣�*�]�����r������+��"��8���${��Sǌ����4��R�E�� z��[G�p��J��5���Ǹ�������IM���u�ƍ�_��4�i�{�v���]5����{��ߎo�.d���J`��X�]�;T�n���Ӱ�Lg����`D1Xh��Fׇ������CV���X[#��a�c0�}�kz���0o�sP(n�G��,��;�v��l�kDې��gʌ�Z���/2��Xn��ב�;��F�k}
_� �j��{`��Lo���x-�|r�_�VvL�[l�2�5qˠ^�F�z>4T\Y:�+�1P�0�t�Ռ�}�s�����W���qG�_�s�o|��ԥdv�V�z��Ӧ6�L�����q�+Z/�6L�Tڟ~�l��Q��!��\>�f�,���fi������>�S�p!VF���Ct�+���&�pj�,��+N���4�?��X��*Vg�>���3�->�t��	��m����Ҳ[q�G��S7�
Z�f�VQ���N-�+A��Ls$��k���[��Я���T�~u�Mo�:�i��!��Ib�ӧ]�=HC~VF]"[�� 0B�z��KM��M^�]I��ey����FuֈvU߬W��i.��)��8�_<����itpgoYD0����|Àv�;����Fb�d��a&(��1l�Z�tSJ�䷛���B��O����1��}{܊bX:m�T�q��^*
��Z�<$T�� �=3*�;�UwO��f�U.G:gy��z=\��c��qB�p��|�]�0mwڅW���T$J����&A���WY~���	���V�/G�}�7(Q�^_Uap����)��TtKݼ��	߭A3���Y���IH!��+��}9�
=��;үH�y��b��/ɨ2��\{�gQ$/��]�-�����<����������&MG8��L�GO���e�[��Q2Q�L�
p[���*1L�0�(��?5nS�ןH�@�ڎ�L�6�3�҉�{l�wk��`P�_T����]�g�B^
�>�\�W)�4���wz��X�g1��'�#O�n�� m5���n�������t����^T-gӵ˞�'���=�9m;�����%w:e����3� լ��3����f������Oq�S��ơ�Zf��I��k7���%�������F���T����u���3���6���;�@�e�)I��Ž�����X!cImpz�#���_��}���ş�+}n"!L���Y��a"�F(G ���-A���~����1,�O%��%P0/���� �A�[��n��SS�2{U�H�;*��l�!:,1	)�c�y'U��>w3�7�+e#L?n6�S3���ۧ��)���z+m+�	�b��)ݢ��1+\�v�.��b%�j��3�׿H�L��G��F�&u�Jiz}�A�dR[sYYK&�0�?����O��:���^�ב�p^yk���`���t�n��h
� �8�_Y ^	_?|�<�h(�w>��/{�}RЁXܴ}��#���2�q�J���*�M�P:�D�g�����E�m���za �n��uo!v��b�MA=N����c%Nm�TM<q 6O��؃�8Z"`��������Xw_X�R�[�S��Y�s>%~�(_�"�u�����)f�D�Ѯ:`��oPFϟ�q�AJzu�~��StXK<%C���kl-V�̇5�i���Y���V=�F��׿7*���tc-����j;\�0+rQ�Vo����m�������Be��K��fΑ5z��(�u�?��Ԕ��e���UD������+�_1��Ge���Q�D���ΰ���|��u��&�5ح��Q�T�2��bԚ��n!��/&^�o[�pU�_/�5`n9|�\E���⩵�?u�*�̃���0~�L�t�;�k�u�L�YJ�q�+B|�݈��	lw�����k97Sc�G��S�B/5�ba��p
z6���-ʦ���}I�X����GD
��~�F=�����9ь����*a5�ʄ�;J^Mז		k�C�p󌿯����ZMG�m��{��U ���feq9+���Ƹ��|��Sq�mI�V��Ζ�N^��Iܛ�!�(u��԰z)�ǫ����5�n-0�A��*Ә��k4ƻ>
tʆ���6>���\)�1`��	�%.}�+��̽(��ϸV&Iݩ�g�����&�KJ�ڻ��4/ �5��	-�`����&�/�'�γ�W�p42�?��.1�оp/ֶ{ٸzP(��qBn}1&K[ן��滞Y�Z��*�&���!f�/�H���h���#�$X�&@�����=b�7��P����/q.&�0�AKGH�GT۟Kd2�r�d*��,��Tf�fk��:�Kq�Pzظ���]�M�05�`���f]I���Γ,�X����AS���8�L�%�{���uw�>7%�2`gy[��k���ᱺ1^|��B�=�@J�-Q�~�ѣ�>S�ƴ�����V���p�,a��o�.��#$��l����N�բF%�*XNnk�n���Z/�[�S�)	���GS*��"��_�N�N�X�U]������1�YjBON7KBL����
,�Pwm�V�(B\���WL�o*�����~v�ʡ�(s*�C29Za�'@� u}���Je�h�W�<AQ��VZC��= !����vy<�֜9k��m]��iO��d��:څK ����}��/КP�X��6MГ�f+��՗ä��Bʳ^�+���)k�0;�׼�p�i�.����S:���h?�j��	Wܽ��j�R�������	Z�yiv�`t�PΕ):PrC��f�jw��t����G������R�BR������r�s8�=�NN*<�j�{sA���~�	Dtl^�DB�z �j��#�\<ܨ��,/jj#�$.;�h��G$M~�EL�(7yBul������aݤ��!�f�R��
��˷�3	��T/�����1���|ׯ@�}��Q.crx�����Nǃq�!!��lh��p��$iEDq�T����\�~���_�q�v���W"R~����_!S
1��D�(�Sn�{H�ӟ�܆���)蚲x��*0�kg�B���j�%���5�`>;#(�� ��E�[GE��}ã�(�GPA��.��T�K�CTPRIi�f�n�k���f(��70�9��}�k�,\�g��������{�"�����	HI;8A��yfa=Щ�Y$ku�6ZN���f:�T�,��^=9׍�ekїM�qBٿj}&�LV��ք�oi�4��{�>t�^i3qo�������E�Z�ߖ�v�ݠe�~�A&~�K�Ӂ"�@�_���g�r.�êY��a������h!%<������J�@��2���ӷ���B��d���T�܁F�8�he/
F@�ad��e�����Ѳ���Y�RtC��B@R8w4RZ&��)�`�l���޲�=���?�[�a���9&����j���K�����5�
�._�K��/����G9:Nbǩd�W��㬯p� �����JC*�v�0�9Csq����-��~@�Q`�C`�"�ʲ��%�K��,�6�=�v*�V"��"�i%�{�"�ŁP
�fA}�S��QhlL��}pLv��xӴ�zݎÅV��,�oQ��k��~;\o�
����o��
�P��K�����l��
�Q:�<n5�&�B���������<|ĕ�4�C?n ˅�i�
���������l_L�"G}5�4�ԠJs�����Ƿ_�3����a��	Q8��J_*��Mp��er|OR�z2���OS�+�6��Y B����:���ҽ*���cX³��*K�qՓ +���>}��]�PI���]c|<����%i ��sCI�r양�rG˘F()+�L�U�f��a�����T�ڊ��k�� ��O(�A��[���e/��o3����s�X�*�^�~��Z���u�d��x����^�����9*K�+��l�k�������wO�5��OV��eZ��D(���8>���?����kۣ~�%c �g2zw{��U0�-��2띴�کP%�h)�.�2[����ݠ��rn��c{��n�5�2�mɤԧN�d�,�z����W !2`�w,�Z�z�],���s���]�T�hu�p{�h��LpI#�y��`�::�B2�5��<w�	��'dg��y���f�>&�:M��+��M�g�Jz����y�+U�X|��|�f7�{cY&�Co0嫥��2Ն���7m��r�L������@���+���`����*2=Y�R�s/��[�\����]y���2�$����%r�\�8�C��{]4�����_��.����Tl��E�?�t��kRT����M9��QT�٠��ց�9l`d}S���3�&)uF~;��f�s棓�8�~�j]ʝ�,r)L������ƞ6���5���ƮR�˫sG��W��P,]m� ��$W̿#B��"���H|�4�l|B��'��>��f7�G�+�S��d�z�+l+v�V��Zb`�i3Υ_����]���_��ת0[���:]��3�~�X�1K�7Ɩ�j���'�e�(��/3�Y��q��J�-Ixٝ�,*�Ƨ�`�$���c+��#�Z'@k�,!�az[,}`KT�E�nXQ����x�-&Ma�Y%���̓Zs�4v���,��̍(rV�5N%gؓY�5M��!ߜڛs��{�q�-ľ|���D%Ax�O�<׿�������w]5qK���q4�eTdW��gʆv�hޱ�����&��$y+m=B�yػ��h�qiFR}Z��xA����5�_� ��9��Y��g}{N���̢��ʊ��i��X�i��pt5rl�In�?x(/@u���:|����!�}�W�[y�Lbg�/Wxk%�w�����̚�,a����-S��.0��tR�]�;��S�\�D�"J�ܩ�Mv��؍�����I$.
���rdؖ�q��$�{�25�b��KG,���r��q+��3��<�fX��^1�L��|�O.�
�mq���J�6�2ލO�SA>E-,��F�-�~|�q����.)P)[ٳz����D!@f����m]���  ��i'`D:z���k�D}��a���prF�h��<����/��|��'�I�+N�DSؽ���Ʒ+�Li���!����۽)<���^'�
%��ɝ�yǎ3��O�P������P�'�Jn�Š���&YvjQ�c+}���T�sp	��:�������6����-yr���8/B����-�0PG){ �C�5fɛl!���+��vګ�j&"��|�����#��K���#Z�y���i�L�W��� ��t�5\�y�i�K����n �j7���� �ѧ�ӧ���ܘ���d�'�x�f��$�P�{S�"�X�#5A"h>@���z�����T��(���R�vv�L)�lٽ�d�$�.k�3.!���(��.`�c���X:{l)%������ӎz2���޲T4�#U#i#"��?:*=,��aj ���G*6��:��51G<S�
Ƴ�7�WI�^vJO���+ը\���9	8JwĿ)���p{������,p�	c��v��j*�,ٷs�M�=�y�5�M=�.��.n�6��ql��-�Oo4Y� \Ĺu�,7[~<z?J�&�� ��
Nh�AJ��\v�̦Z<�;�8���]Ł��@�[ۻ�
����ӓ�i�\���1�ffi䡻��`�(7�,�OD��l��썹� �v&k���L��g�h>�3z�����U�#K���;�B�W	�5�&��Q�1��S54��,�3<Ogx>��!�6�m�?�=�L$��鶔5>{�Ǝv��(/f;�b�Ł�+�xA�q�/Td}*�ZH|�<X�	?�a>�z��N�c��~q��%O����&C�0^Q�N8�	
td!������PH5N&���q&��ᏪFU	�&�XS�jZj�H�ko����.}&I*���!MjQح	y�:��&�a`�l�,�1��G���d���4S1,,TJ��	�*E!����&�J�"�E�NF����P�S��%	5��7�v�Ŋ"ڢg����6�ǡ�y��˒_Y�t-����6ˣ˨�(>�pE��G�7Cw�-�����[b�*ܧG���3����;>%�MA�(z�I��/�E��P��|qP�}=�I�9��ҥx�!�X�[U�On��ѭz�gK{j�P��U��Ðwg}�qɝ>:�Ď�8{}Nx��N
��� F8�8�ꚨ��(=�Q��u�$� ���+���~YG�����#���ߵ�w8`�4��5SҒ���c��׾���u�"MJ�0����!�.�nȇ� �Y�^1�/�G��y��^��8���w#��ӹ��T�;��ϙ���dE﯌���ȅs
XTНB�u�l���/dq�zi����فI@��͛O-)�Px�W�P�4��[�K-��i�?7��_�TUBp\��N ����$��(>)]��m�0]%�,;���SE�R�Y$�G����T8u�'��f��(�fĐ��mGL�5�01��}Z��f/jxw^zȼ�$@�|x!:>�č!�f�O�z*�L���3�q��N�!sy �*z�	{�Y#͡:�u����<�,k�+�>kmԭ��7��2/�#������.�s#ObA�6��o@�.,�E{��1[ �f�YXO��ɖ֨��Aw��Ŭ�#<p���W�R�s����A�9�قKL,��NE .!�l��w@x抭����Ԟ�(>r��s �爙�� ��8q����\9j#�{6͚���2�z XZ�斛���_�L��M x(���xo��@������W6�Tp�6K�Iܢ۟��Z�BJi0Ӆ�ղ��"tֺ:��<�ϓ81�?������"3�ݚ��uKCeMI��*����N������>YZ�2V�?����N�%� <����VO��)��N	�7��S���p3�����q�L<s���G��r����^���`Y����|��i��yX|��C���(P���O�|�\�Ê:6��ѭ$v���e��6H(�d2~�u�Bz[,��QU� �B
��*$�a���n?̷=�0�%; �f��74�E��d8@�Lm��}�N?��k.xRT�HsX:��1/^�XR.�mz�.C����;"G?�E�Nx�C��Y@b-�%�p��oŐ����a3T�J��� `�!^(�\����½��Ul�����mȱB��q6�n���P��X:�	���B�U;�/F� ;f�*�c��}޺��𱒜�5d���8���8����&;)�CY/���q ���
~oki#��8�X_����M��F5z�j��3y��g���{��]QU5���kM��d�Z���m��?B; �@���={�8|�"G3B	&�\�_�q9	�ڧ룸'�X�^J_�����U>��7+8E9�Zk�/��>b6H�m�]��=G�M���O�z��JӔ/��=��7��`�}13�ؖ�*<���0h._֜�"D4��H�O�병<�-+ ��[�s��Q�N ,L~j�2[�"��58�M4G�׈���Bl��>%���ӭc�^�_J'rd��ۭ����6jQ��H6���G��,J����`���fg��F<��ī��Z�R���&�+�\���&�9�
j����<,I��s�o��N������ڭ�(|����޽
�������~���Q�Y<_��պPb��h ���ص Gzh�Tqf�\�)��\��a!�n����G:�h��守iD��������Z(��(��*z/����:�?u"5�:���$'ݓM�p��k��UN�w��>e�H̀��r2,���0���P�vl�]C�}��vyB�iz����`/or&�7[�y:hwS�y�Ez!*�\N�dU�ܗ�o^&��,��~5G�ァ�ݽ���Bi��i�Ç���M�ʞ��|�Օ�����JS���}R,�Te,v*^�R�D�a��^V/������֥I����+s!:*ʳ�-\�3@I�6Ә��ЍzvwO��>]z"�y���{��z��h��:w�na�S橣��x��Jck��D�S�x���d�����+}U�Sq(��3����R�6�q)liE/����p�VZcܺU�OaǑX?�Z���k� j�2�08U&0���j�O �p�*��}p��̣Q����Fk���W-2O@�H<3}����Zޖ��{��O�),V^���wy�j���Îp f8MPVv%K(�E�2�tI�`��c��I�����p�Hdn�#�ي����4k@kN��z28'����Ie£��� ���Zah��I ������=�}�i�.�� δZq��T�E�i���iO�L�t.�h�H��eqz)C�l�.��t`n:L��X*�TE֙aH�8��M�*ѡmi��ӕŅ̷��jd��@����\��D�%S�4�ſ�z�����CR�����$�O�.<}�q�Q���8�K��<��}[��QC���d��\�80Z=�F]��G/#;�׾�ح�8�30.0������v�'��3�2n�t��V����+�p��.'P�Acf��DPrr�+2�D��'��z�!����S��.vKRBpyHn���:U���-D�A���wu�h�i�n]V�|���z���A1���WZs�������o6��ѐg�"|���.��jY����B�A�y�~��N���ϱ�CEs��~"�@y��?��L%��\��T��*��w,�f�D��)J
����� �<��
S.�M��85�:-�ХD�7�9��R��W�� �w����L��p��I�}�
+Vחɫ�g�b��נ!2ܒ~uw�bv[�bG���qN����s~i�W��jD���G���_��ò@�b�~F��}����r�ۧ=�#:�%"׍�g��L'�����c��b�u��x�7�_�
�47�PIZ~�]�`�*��R�co��P�*b�wO4����a���#�)Mv���;�k{�fzU�k˜�ᬭ���!�|�S��������f�v��c���h(C��������j���Җ�����퇿n� �C�-Ȼ�_�k�hsŷ�b��#�U)��-Aq0� ɽA�#J}�1r���=���@�u��)2F|����h}'�/{��)�_������Hb�a� ���X���� �]���d��r���I.S��1`>��r���*��^�Px�ƚT����| )3;�/��O�N��+����*홑C%L�h�|�z���ik��<�W����r�Z^�=氁|H���R��a���?���~G��C$�_ߥ�Q����\�9s�%ǅ�Z3�~S0eUG��۹//`�[�������E�ݯ��|��S�#|v���iKS '$Ee�A��h�K�#�-��!.�C��¯�t���E�,?���=�W4��>��R
����RI�b����R�epB���K��)�����Z�w ���
S�-��l��N�,�
ue�難��20~���a�e�`���$�^"L���T���������a @��

�ឩ�w�hd���M������!/���s�?^S��P08��\[��r���Z�}߼M��|
����q���RdnY"�[q@��q��T�������B�Ru9��x���J��y��v ��/v���ԖP�\�B��� �t���Tyj�b~Lw~ORm��2�z<ų��e$��� � iW��c��I�V6��A���Y�R�4��%,�A�Χ��6�Zs�~���K,y�}�]+�a��Y�& �̷Z?4�W����$h�x���N��!wG�c�Ɓ�H{C}eT%�}��R���n�I�[,α�9�<��K0�@Si@\||WC�i�s��d���j��Sa��E,	�ʼ��v�'���Y��}yq�>�M!d+y#P@7��s��T���%���X<V3"��z����4�A�P<��q-����o�6)����>�|��|�ф<������їp���b�	��-a4�SX)�}-晢�(t���m��Ed�P4�	9f���eK(|RL����bĔ���F�]W�ࢧ;�}#�-a���	ҊoŘOwNލsh�?4j:V̟Pb��`��P�y�+c�b���H[��'��}�\���NKi�4)��F~�$����z�̟'Š��c���l�{�����:=�p���N;q���,5��0��p�OL� �L�y��������!%v3����kSV�g�I{��ʰ	���u-N�3���j,��O�M�,����9�$�X2q��+���h���9�Z���l�ՠ�{W�Cb�\?Lw���nd��!_����ً�ڻ�d�.���G���X��Cf���aӝ���k����S=W�y2<��7�J����vcG=z�������Ԛ�Q1���%`����c+}{~7�6=��Ge��+��_��o�(�r�rS̰!�y�6�����b�,c�p���|��«�ˀ;xh�щ���Y�6Ou�E�-�ͽ��(�� �����:X�4��%���i_�|r$���7�Q����D�T��6jnK�*S�Z��;݊��= �y�֯�X�+w�ͻ �#��={p/cz5�oXiN��@����_��d�D~=*�=�%����ɩ	.9$HK��}��/֤�l\�5`lǪ��Q�9jڏ�f+CrP~3�o�]bsQ��y\�gQ�ف6�5��I#Ji��cY�VC�ʱ�Z��Z�lFӜ� \kuc�\�����wT�n]�׼�z�W2�T=���ϵ=e�؈�F�-�`�S�[�L�.w8g4:���<����O���ܴ�0,�Q��D'�fB)�e0_��*EEEB����9�YSmg��c@���xQ������y��*�D�����P��&$_����L���L!�J\<�B,/����]1W�Co����2���nT��C!'ޜE��b��-��b�U)�%�.ӌ���)1�h�FR�~M�y��(�b9-S^�v��O�A��_v�T	������{�2�l#5�����B���˓=�^�丌���Z@��S_˥�eg�o���_}�-p����|$�>����<I�K�7���k�he��&_��{�!А�Y�xa�iU��2 wC��;b>�r�s����Le��-��ݓ�y�(�_�e�� e�L-�TnH�����z�ד���
aE�,��k��n""�FA
̓p-���?1�_��(�9�r1w��i� W�Q�`Z�Į]s� ��E���\� *)�B5 ���C�h.�$����l�\�4O������E�EI�Eb���8͹'=�'HE����"Z&3�&�ёbS !@n/�@���t�
J,~���f- ����u�� �z��f@ڗ�nsqg�c�2��� s�������+��TtM]CE��������a�λkFS;j\R�+�HIW���>�%Y�b!�m������z�M,�c�^��N3��B(h���ʹQ�Y���~s/S�&�S�=Uh[�I;z� we�g�ف{>�ҲO(.��T�*u{����ϙ�yj�Y��2`�B�>�&�R�ck׶��sX�TliA E�P���S}Z(
8��4砄����<-�c_�|<Y��%����G��T]��؅uǡgpd��ݧU�E�wjc��'�ι����#a�<��X�'�$XN�&�4�8�[� �X���n#������rEm�_[I���3�t"KU@�6R��]������n�HI�8�0`�|�q6~.��[�8�O���VF�c�ae�RT2�jh�7���\�0��uf̀���e�u7�ϗ��A�t���ւ�+�pR$�ʥĐ^��A��9��t���\�{�2�h�G�Luv��2�/^ty=߲l�'!X:������׊���H�U%oW.�n�=Г<X��nUQ(��*^tٴ��J�༼��Fe��W�08ja�y��O�K.-�;����s�N�� ��Ԯm�?Z��}�2���A���<u_�su�0XxH/@P�nZn��ӥ<t��{>Hr|W�@�0��nH�nxOo���>����(�����TwiƗl\��O2���֕m�B���gX�:w��l��D�|��D�zd�I�4�V���&���H��O�$�yZ^<Bo(���g�����\��@ة�=����p�J��O�T��2ܪ��V����N���E�RY �/�ٿ ;;�fou�^�z���bkK��N25;;�	�X3�U���#�5�+`ܱ5��+�W���F
�7��Q�Zۘ���7ߕ�Yb��N>Nt;�\�r�u��HL�zU\��,�<f�@0��=Y�δ�r�I��|,���)��L �8�9� ��⤰�����1�Fw�"��I���5ϔ�P�-��K6�T�u��X79���&��U��U3�O�VcPn�ٟ�۟�@��w�VQ�;���sz�XX�R�-�F�5;ީ��t�_��C���nF��/��|ѕ�=ةe�^�w�D������?O Ǳ�/W���%��!�ð��~ �o8����:[c.=�}KG����h<̈���t^Fq�c�����"w�c�[KY��/����������s�'�iD=����Sy�Q^9�n2M��сJ���������m����>S�.QZsY	����,G��֊�|�;b�=]-���T�b[�0��0�RX�ʰ�A��ی��޾w����\%ɲ�')���7�
��@�&-/����6O���Kv H�xR��o�\S�1ބJk��}��B^�L��Y�Th�騰�'�'�dMi���Wʐ(u��&�$���JS�fJ�ҝG�����SYLe� �T[��s0t��C4a��vw_�m��!˂��W �`Gi%7�2dQl����ԉ$����@���Cko�z�șy�s����W�b��~��;n��3��� �ߥ����L��ô���X�!�I%�3�8{�1]M��.�|C��O�@~e�B��I0����ed`��Ȟ)�b���88����QӼ��~�QN��n5�ޝ�ThA�(RV�,��^�qP���W���R'?58LS V��"��@���Hgb�O'M��RȠ��+�yY����:k�Ļ�~js����Ȧ�su�;�v�ف�l�3<�}�yi���*�:�*b�i�d���p:�ȷ�'��$���U;�|����T64LC@�g�8{5�=_��h�E/�JB�u�������=����G>V�j"}Z�.xG`oD�-m+
t$#���������S�>��>y1����dLR��|>���<�#T���h�H �	�����~�ӧ蕈�2��%�j��/3Ŝ����0�yŪ٪�c��4'1۷�n�61*�,��i��c8�A"�v��p�����2���EW�
���G��bB��C�;�����	: ��Ju�����x���G��FA"��i�z��wN��zNN�g�fo��
���-|U����6�g��Xr�⃮qCc����~r]��i��<p���<� Ή��:��S��nټ�o�6 ArE�� ��I�M�?Dh>�T\f�S���)9!Y\D#ra��dy����|o�#�R�:�Rj�3q�E�	ъ(�gY�BIW��!!\y�	�PV�6���6���MZ���Y�R�J7$eb�Kx�4�q)b0tK�bc�d6]9�{n�g�ơRG���W�t��/���IL4����I�3�lf����W@��ϴ9�GWkx<�I�����:k`��0��О�{�2���m�W������P��� 5��>Ԙ�;��SMa�u���O���0��޴�}xݶ�� ˺u����[��L��q����$�|���71bc�Ů��x��x�#���n��O�8֛`�?y����^Z�����L�$u������q������7|_����\�Ƣ��(�I����+�~��R�6#k.�s���qC����>�F�ܬ�g�F�G{�;?�,�v"�	9hdÖ+@O@l�U!�R�\�>�7���c��J�}[Ǜ��{����;�Иj�P���[̲��I�.�!  hLԒM�r�)�Ch�O��PȋN\H�i���l�T�qF�8��+~����L+c�����/+|z�
D@�U�P"�`�=~X�4�(�)���r5�}� j�:��*=��U����QI�>���G�~��
��b�Ο�)`o�ħ�[�μ_����p�LC�36��N�h��58�(�x�ڕ5�peq�ݪ5v}�4 0��^=0)�F])5���絿��db��������+��u��Qx��Vf)~W��4#U0F��te�p�J:�6��f�K�Tf�H�;�\�����b-�b�6�K�#� ��nF,���٪�p�m{[�e ��q��s-�M�^#�Q����g��ϧj�n�U?>5��Rl��	�4FO�ᵵʪ��M���KŢ�L��^�2]�T'ya��9�,`}'��8���E�3w<���T���W�V8��rXG� ��/Іve�Sz*��5�N�x���q��(�N�*{��Ry��M�%	�{�E����P�78�����G.C�r�g��(�{�	TH��
`���]����{̕U���5D
��DRr"�+Dz����w"��?��5�G��Gk�Q���u}���^��}UX�����q���R;�iI��9�xhB�D�&4��'G�EG�*�'��N��L��'�+���;BdR�D**Gu8���EHN��]���?��}|3��x��Q���I$f8�V�	���	�}���x9��a�����q�Mh�E���"�f�钔*��Y����
݅=ۢ_S���):wL�֪���ejD�~�d{��~t��������l�)p���li��Z՛����-�T�3�_�	d'`��R�˞J3����I)|�-�c�I����������/R�q�s�����B����N�Y*�N��_O�b�������?�I�~�1RY��� ����m`��g,4g��}�0t�謙}R���n��]sYb��n�,���CD�H�r0_������ɛO��]��B��u3���k�s��s���3����Ƚ����P	����Z$�T�Nі���T-����C�L�#Ϭh�G:L2�$�b@=CJ�}�v���V��˜��Ψ��,G��?��pv	h�����߷s)l8�z̢��P��y|��~74�-�k�e|G;[���W�x��z��KGC?fQ�"r2�
�R�n�-�R�m���f �����= T�|=R��%黅Gԉ�b�֊H,�1���ق4�������sJ�",7�uDh���j;áZ<�B�@�3�W�#M�h{P�E+� �V�l�N$1���,ӰNq�m��A��x0��;WY5��{��ʨ"����Ș�L�DP���U�s���J�(+�PV�=�C�b���˯<yX-��-ĘuKz��te.�((�&>���{)��K{1Io{#�0,S޲h��� d�o'�� ���$�ƀm`�����!�'F��;I� +Ņ��~nS�bZ�5��(�ڟ�.j�Q����?g�	V�ϫ�[p����"�3��_����"���v�J0�]��Q�w�t���9	�W%v��#�(�/Ei&�q��)�i����0Dȧ������aO�3�8���۲M���[�r�;�������L��<�|�4ϧ�Y�}I�jօ���Z���Ή�� ɽ��+��UI=mͻ�o�^���������l�r�g������\�ԅ�ۜ�L�S�0Y�SIl;� ��O=�p�T�vǞT���rph��OAf^B��4l�Ot�t�?L�M�Wa�2�"�Z+`�a��}���4����v:8�cA3�����V_��gfg��2�:���"�m��qꙎ/U�� �6g�I�ڏ��锇ʿ���$�j�T�vntt�v�3��:D�5��-�XI��\I���C��E��N��B2���%�]!�J1�rN�슥mb�%�~I���0�Y?Q4mm�Z�]�^�fbz�d��F�ٷN*��.�N����]i�h:74\џ��}���g�6�Pa����;��1;/��LR30���x
�?�T�E k� h),z4L��Zǵ���=/?^k�I��>�;٢Ƞ(�f`h��
�A�u�2K̆�K�DEEÞP��P�3\'h]�� ?l��>�μK4��[�z<�o���V��X=�|q��z�h���������g��xR��q����n�_-���E��q}��4�2#�Z�#��eK{=�h��=@|Ɇ�Q�S|�P��|�\T�u�����i-�vp(�n�	�gRcȭzfw�{؟+�-^�E��kʹ�||���8ǉsv�e���|��{��9Q�f�� ��I}���%��Uʃ|�s-���l1�p���w_�d䶱��8���F`�K�AO�u�ΰ�?y#��ܜ�`���,ex��h���hkn�� 距�JdK~�2��t_����|Y�
l��|��v��!!���������?�3<l�?�!a6D4��&x'DF0���Y$�wp0=-�9S2C�������ɫWihlD��̭M�����x�.W�԰�<,Gon҇4�����cn>�JN�#�ȶ��O^�I��W����
"V�'r�'�"�,y?@e?	)����XU�D%YŸ�Qp�ؓܐ6�H��qJ�_��l��[1t�:�ͼ�+;�lt�v�v\! ��M����!�F	cǽ��2t���`���8�����Y��r#�/w�Ō���q��Ź,Gڇ���j��	�F�/��V����;�/�ˀ�|�Ds {O���-@��h㮖��k�xR��R3�r~��W�.I�4���{��i�'�=�iX�`Z���=��LUT�Hc.�:{A�.������ׄ�l���^�U�r����W�7�M��2�J��z/|YZ��F��h4h��
�\�2�GU��V�j�"RRRi,,,2<�Č���	lw���;� L�v�>鈑�H
����?�z4��h��֘�d ��b���L������&�m�3f>-)?�*��٠�W��ܜ����ν�Y`5G�K�z�xC2�-J�nE�OM�a��5adj�е�w��7�Ae����)���|�X-^/2�}�П}�QV�G�(B���q�b��6޿�f��{moC�����]���R�ߧ�!�V��R��_yfcl>��,S��}��g�x�D"-��8����l.����x�귆�B�\���.�<�}����/�&�T���t
pg����LLL����#�H�q[H���.z���gT�:�ҥ�1
��]kW �"~WRb��}�9_��3S�����.�Wy^�劖�����Y��y��ҥ���n$�U����J�6ЈQQQD�;+**��{�Z$�������
��#�����!g�)�ħo��%���$麂�Z:�hO�÷:^V��H"�Vu� Ӕ��5[�R�����@]��`5"`�!ӻ�X���n�8�4����?[����8��L5���V��n����������%f����t�#�AL(^7�C!pk�sQ��c�z������S'�"��^�FD��塎���W?�.��c�q�p��{�o�׮Sy���i�@x�*ig.��GOV�7�E^�Nƕ~�&�Q��)�p�q��������T��&777�"4|�J�'65X���j?ʻH{���Y�e�xWkM�n�����_�p� $����!�`0��,���}gº.0��kO�V	��̱�-tV��$�[/*�J4F��Y�ս-J0&��M�i�p\���+��Jy���! +�:����P�T:r9-�^�l0���ɖG������;���׶��*$W��H��qwX�E�1Ͽ��J��1��X�j��K�{�(-�ݹ��?���C��ф���gJ��� �UN��_���lsqh^
yJ#tC=5D.}��3BZiʽ9���������3�r��"��^Z"�F 
��.fH9�*A�-���މ�x,��g��Vjv <D��4�������*=�'��;蜼63u���EIFn�����W_����`oK椧AM��}���h�x��C��g��V-ti��.P�8[����B �'TUU�������X��>`ͧp��C��!��F[�$����?�R)Ӧ��6U*:��:�ӧ[9e�<Y������.�]����%�t�k���`bN����]B���O��E��/�Y�Z���L�S�\�~����r�lÐa|,8�Q���?��z�N�=�3F����Uɚ�yMS�&0��
0�(
��_�~��1��*:c��4�62&�4	eM�B�)��7��S�iqd
i�R�������:�yԹS�d}��sr���m�bP�'6zed�1]�I4_��vRTS#��q��%w`��|$/�_BQ�7����gHV�8��f`��Y�!���I �t�{*�'���iB���"�'M���g:K}q�l̷�ׁT : �G��e;˕��Y������!�вWR3^�_��|���=k�/-�z ��ے�����2g[|�{<���kk;�����&����&�z߼/X5�;ԩƆ�=����n���615�i-�/]�Ѝ�.M��jc�#��}w5��:�������'�T�_�&��v]4�:��L�;�`�̤�O��Zo�nL�� #��|�>95!�FN�Lԡ����6n�Wv2�u���1���C���y0���m�,�V&�P�����z����n\*L*.�\��>388�W���e��{{���T[� E�q�m!�R���ZqQ�a��,����j�~��e����7�s�7�w�@w&[|��r5$~��q Y�}�E���e���QaF�ncUNV٥4\A�Ɩ��u�0�-""bUO�����Jz�w�Η�6\���Б�N]���շ�u߿��erV�" �#%B�Lgw��0��r��W=����{%R\����^��O)$0.d�7�:��l�-RNA!�����I�ko{zz���4���f����#��(�J��� Tt�GƄ5F��}�	��Gcyi�?��Vio��Z���
��9Y�����4��yGi@�7&,�K=4�};=��ߵWm"M'����Qh9�D���c<���u�����1Wܑ�m2(<~��Qz���M5�$%$��i������oՂ�̵�K�i 	J�=j�����A�8�*4l$�����@�e�x�0~�1߉z��#"Ybb+׵�xP�����	�ZX��Ht�J*y�@$��z�t^
�mZ��xA  �!����J*Z)#c� �iX��^-��s��`�]D��������z�]�44��ñ��Cn��I�9��Վ���^ /����a�o��`�l�z��6)H�/?���f����z'-�o$�ɭ���R#��
1�rphz�����L����g��7�f~�% ��u����X��������I(�[��.�f\��wƶ�}}}n�;ȝ#�<-����Qy��РZl��J�ų=:�z�E��Lrb�Y�������Ttt(!��;g^x�ޟ����HyFV<C�K�b���%!Lw�D���s�Ѵ�r^P� �T�޽�!`�ehx�c�/���an��i��GNS�O���Ó=,o�dO	귄:�7!t�.��&D�֣j$���y���J��Ptp�l�yyw[Z[	#q���6��[���w��!X],��Ȏ/R<�,r�j:L�S2�V��m���<�������N�!�~��WPP �;444����Y�s�F�^���~������t��KJ��!jg���;GHS��V(��o\]���P��5���Wg��KKgdg�����̯C�	�%���*WF(�6���ޟU̒TS���q]t��Z�+,�/tFq2�H~|߂��q����5��񇌁��R8Q�cz�S����v5
���)��xy���:����1�0|͢�&�������fm1��a�!	ߥ�
@y�V;����^�ם��@���
��溍$��C8�4�K|]�BM\���o` |����Ռ�Q��EC?�yϛ�-;�F� SRR�@0EA����L�����2��p�Êi%?��n�!���!��}5%Bx��b�����ɷT�O��d��������z��F+8�І�Q�aaaY��؇��X�|�_1�c``�.��d�r��^��.P8�%��������Ei���|A
bLղOKs5�� �8Z�\�F�� �
��?d�Ks�7�,tl4���]�I��7�ފn�_� "`��w�̓�xGlO�Xh9�-D���6��uK�Է�k;쬤�4Z�l��k$' N��lqq�h�6��Ҭ����	M�!��65�����(�L[����㝩����֏D�xPa����:�\N;�05���GI�f��V�tyF��\�95�#�8���@�K��>�s��+�;�����)�I��d�rs�cKV����Z����a^.��m�r%�B+�a�j�sii�[�����W �6���.2���=���l��RaIq"��;�G�O��x~�58�d+"�%�U��? hM�M���볝A&������y���+r��o�O��f-˺��P���UD��Fo��k�=����p,3s��Wܨ���˳���W�lI��
��0-�U�p~�8i�Lg||�P}���恣��1pq���Z}s�$��[Z[g�wS���%��;+��s�w�-�;bڥ��R�N7�,}�Y�X�:v���8�����ӹs�׏�+�����,���箋h�1Z���Q��'im�y�t�uZ��C��qCI'��=<&������-��*i��4�gҰf�L#�����@B�����ўX$����R��ܷc�߾47�3{�I��u5{r��AߟS��ZiIC����TEho7����q����_��kw�i)��N�f�������k��W}��HQ��R��⥉tiB(�	=� �NP�R���AzQ ��[$�WCI��?'��_�b)�0sΞ]�g�=3.=�Qt�!dwx-����P��{r5��"��j�|�AX����Yj�������kV���k�e�),X_`�Z4Ғ��ѐ��t���ĝ�`�^�����ƾ	V�����_��2��j��>:
��Ž;1�6���V=�\�ճ�G+� �5a�e��Y]]]k�������c���1�7 E��0��*@�gK�e�"h���_�
G�4�4�
�����Wbz+����P���:ry�9�������7u_n�f�	�H�L"���v-������1(((�S3Lz�� ~�<�c��oXj�������r����yS�|�=f�*�����k���/�l��7�9�W��^(Wc�&�U��#�+�����`o7!��46�̵��w}�����pU���L������xP���*-���!��,�%���`U�C[�v�~�p�"��<��^s��3%���[PO8�^�{٩����/��<�ޟ^�k�Ř�z��S�f_�����]oy{\lz8�/:�:-]zQ�|}:55!T���ƖY�Gy�A�=�C��+�ڔ�i�Q��	�lO̮����M�m��>�lK�_�P�Y��+�J��5�܂���3N���GX�h�)o����<C#҅�X����b�go��˗!AɖC��ۛ5��嗩g��uI�}�x�����YO��a�L�7�4*�4�LA⿂�7�����,�`f_�PW�ќ�b�����2�OF�>��- Z_KI�d�>9�a�j���H}y��!$���+O�0���N��A�۲��0�p42A,WVnoM�+-��зρ¨-�q��9�d�����M9`��-�����
O��o/Pt�F^���m圣ߴLX�52�,��e�k���Z��:z.F�iatA�4�z �Sz*��?��r�]�)���@�Ԟ�~���ߣ�m��%�����ޮ����f�/; �#��e�������2�a���o�^{x,��΅<P�n��a{��~���&�\P7�������H������)8�*�LsJ�鱺S�~YsH���K�k�!1uw�i��n�ѵS��_𳷺NgU-9����AMAM e��U]ӥO�Ԓ���P[���V�����M��N3?ۉ���>}��*+ua���+y�ֶ���h����kc��nY�Fvn�f�-�Llf��+�7�����^� ��v�����_:�p���bO�!|"oG���t���{�M�C'�qg�-�p�m��kB.�}�u�����</�R�,s��0�o��T%�� /Z1���L��VJ�!�`u1W���U���`Y�b��]`�_.�a[��o����5# Ă��	�G�bw��.C�6��8L��MFM�y��&&� �TH-�h�ͽ*&��!��ÙL͢������Y�n��:�u}�ׄ��RZ�4�, "�u,T�55��ĆR������_Ň[�h����9Q�C�\�wP�w�c������:<����|�t������B�����[��� �N�_������c����K��=STYfi׭�X��jv:�z�r)M:���tz�!��lU�A�÷����.[�v���e��k���84�0lU�0��穝ƴ���?d�A��
�tH`�(�_����튒4�I��k�� :rb�ѷ�ǽY�H�L� ��e&����|d!��.
�p���J�ysWˮ��PY��Px���P/���Kq_n��~3@n��~N��pM6�#+g{�[ʝ�%kS�+^�t'�4F*�?4��1ʠ)�w�c����!:��� �yI�0LA� �x�K�Q\�.����Т��b%��������p�6y�`v_�R�ߦs����V�5;D�,'t��]! ��FV��D5���p�0�/4����fQ���+�@��M�A�
�[�x�iS��2ɾл�RQ��(zѱ}LD���D�Cs����� ϩ�mhg1����T���hy�׋�L`��_n�k�Y�0����S�k��e�����:K��?��4珔$�F5;0�/���2��PG2�L�ݓJ�����*?����dz����cA��ThX�R7�VD\\���锝��R�ؿ��N��7�Z4C��p��W���j����Y>`��;�{GEE�i�-��݋� ����6ճt��~�~��l�ĩ�[o���`57dr)X�5��2���� �!��J�܍����]�C�$�����iW�����q�^���zp��co�e�(������*q�R1g'M��+v�ۊ��3|����yNj�^���U�������M��\ܖ��i���޻��+!�?�b�ʰ�����
�e�T��0������P7U�PԀXT�����N�q�{�a��EipL������)��m�̎�����	��0��'��PN�}�e�nxBk���29���Ė������o�SH�++������N��E��aEĦW�Z-�sS_N4\,)��}��=J&��U�:f�RGE����q &��.�q��bZZ>�5�v���Y�!Q��V�t����M耢õ�� ;9�����E4�
�blY�~a����5Y��<VO��[�c۴!_���,��!�Mf]�-	<���7lM�T�O�67 �RU��)CrT�7{�1R�#r��B *�����d�:��Ӓx�rv��A��x�n�����ܱ)�	'�V�$��*p�2B﵋;w[(�
�� h�g�d��篘��#���
~�X�Qp:����i�%N\n������]yꂥ�+���f��<!g	?��_\�*�_��8�~4Q��4#9���Ju橇-����>h�PI�Z�Xi��M/��"Z�]�0a��Z)WU�n^�?��|�k?�"����Ȍ8=������_��C�F"	��ڪ����~pLx�zu^Ҁ�ia��o��s�Y�,e�u��5_��FDc����h�2d�����b����U����'$$��]��De�wi�A'��a	���,W�UGZ
]�� l�@q��[���H�6�j�]sEkUS��Y��*2,��a.W%�����}W�0=}��:*����P�EN����y]���r���an��K&��DG����zZ��uſ� 7V���+��k�q��a��&��l&��,rw�\�e�?��?e�-KDe�r	0v/�ey����ݩp&��+T��K
��	��>��<
��� Z/�����:t`^�!�c'v���+��a��Z�����a"���g�T�
A+���5�U��� 3�;���ȗ�]yz�+D`Հ�|��{�l�1J 7�����U-�hgH;60�\s=�ͫ�o�Ǝ7X�39�},M+��P������E������ڛ�6����K�a��J��+����]��a#�/�ve�@�X�R�%�v�����K�L���^�I�����f"f�?��Z�1�M��sHc�>X��w~7� �������Y^�,]�:���0$�ɋk�K���<셦U��U���r������k�ʉU�O�ʕ��y�tT���F��O��}s�ln���駖�}����Y�n����\a���L��7��\��(��������xC"�ߜ����	��2ߚ.f����S_֍�s\<����\|�� ��s��(	l���8u=�No��wb����T����D�Vk�[P�sMm���9��v&�� r�}��N���H��%_Q^��x�H��$�r�|� |�j���4 7���'��P�ng�e�<0�m��;�$л _+J��t�=z{G�r%�W}�h�5=�~�v�:�Q0�t���چ�2>��|	y��'�ז� �xd<1��^Gf��㺟zT��ps΋���4�]�[�F�$/�t��Yk�Yn2zp�������ad��/�n�~���S�NKƬ�zz#7��d���
�O��1��b��,ru�H�	�����Lb@��-�8fZwK��Z����7����䥝�F/�cW�%i�ZP9�O���'��dV<2�v`ș�e�a�@hC�qX�U*+�Ž�� T�U�����=����fM[m�G����r�:w,{r�yM8�N&>5E �$�ڡ�Tף������0��mVQ��:�@J�af��碑��<]��c��S�I�zCe�W�^��^bl��E�*-n��66���0�w>�iS�����n�O�2�l�ܬ�����jQ�f��3�T�i�A�cD|�,��AWx#���t#��r`�I�b�w[`4�;��J��������KG�(&6Z���f�c８i�K�#Lؕ
~$ ��i�wa��ûK? ˑ.h��5r�T�# �h�nF�s�2\EUG]_�ү��������^a::�U֛G�v��;�#b-�ӑl�n1q.�ހ�]°1�۝=�Ym|�J���B��!���A�$ک�~������ݾ6��K{4Ӥv���4\nE��9��1���-}JV�!�H���0�b>=v3u"�[�DU9��G����߭�k:�^�G���e�
�U~��0�b~Zn�?}-����:.�32�,i�	�F����������+�-��� 3�m�e�R�>+A~�'IL�X 4OL��!Y������/%��]���3+b����TS����&S4G�]ec��E�$�6Ǭ`�<��6l�+����Y�ܺ���u�D=>��3��G@�����\�� ntc���9����K!D+lp{�M.�Bd�ڕT��]��CƼ��e�x�������4�n��PZ��*�JZ(�T�X��U��LF���[Qn��noo����a��Ҍ�әO\~7������\:w���~$�9-�)n���b.2A�U��i�6����~\x�dJX|��h�����O��r�xC�p�m�`4�g����;W0�G�֮2����}}��㉭�� ݅#7�  ����$�;YR�y��ҫ���Q5��oH�C����R�z�J� ��"A��5�o
�9�� �kk�@'ehఠMh��������=�@�����eU�~}�۪�h��z�y�X��G��U5뷭O@����~�����,�c��s��k��/����
��/�c�i(��
pPWR����zMO�:] iOw,�ۣ!�ܱ�.K���k�A�ځg9�J4ɋ�*�?C�	��c�g��:��6��(XE&���8l~@�!gF� c.S�o�_>|BU3w�w��k�9�(ɡ��*X\�)5�� 6��ѩ�#JJJ05����>}�"��.���0KW;��-�Gm,� S�-{�Hi��~��ӑ� �h��*J��|��,+��+�B��z��q�?�g7n\·0L�?5����-��=�p�}v�m%��7����~u:Z��J,��)�w���eAN�-�x���[�+DFGGZ���埍�һ8����n�{�}����t��S����|�=@�i����K�v�4������-�k�h�.���%�ɽ�}G]��J3��4 �-�g��5!f����v/�i�@> 7�E����e�vs��!6�?���s?x�,�W�}(D]�d|��@���nȭ�ʹ��\I�($LR�z�3��
�q��D欿��23�J�`���ڡ?%<��H�d��6�i� �r�*a��o�*.U@j�� R S�(���%�FC��a��Csꦰ�G���4fOXp��xl�~�K���3�K\��<� �Y�ʖ,�:�ƶ%����u%?�z�Ԏ�]'�@�P�!}]3)��ߩH�s�kcAY���<��	L$f:qqu
��F��3��_K��-$;�3�"w�����~oP����^� y6��ϲ|>)5�}����nʚ@�(���+��pF�D-#�]Ẋa��,r"�"Y,��I�0G�����%���ՃmHy�n)�i�G�l;@6�-�(��(�n����X���#n<O<&%U�=�RX0��ǄΠ��2 gU��&畠h�u{ �˖����2���Jl�Y��̘L=tK�	���C���w�6�&w������U!�z�_�??x?v�Q�>*L±�6�X�	�yuE�;%1����G��&6h.m�����#���P��uF��lm���h-�=Wr��dZ�l��(��HN�)��9	-WçW�P+��Z�n'+�8�)�:u�Ss-�S�G�J\�w�7�K��nў��s%�Œ�����Ɍ��~�7n21�^_��3�N|��炃��e�Lԝ��hz'd1?�gØ����G��'�>;�([�&6���]_ǔl���$���םb)#���$�~iYvy'�����0mĲ^��K�(u��������Hi���)�T ӇP�X3�X�^��'w5��G�y��r��e|��qg�0j�(w9Y�+�0���c���z�U9�{�E!V!Й�Y,�`w��j����O:4��1\e�� ���9�&[��4�vxt��)#X��;N���0a��
�� ��]s	)|����c�
�#ŀ����9j7���R\\tH�@���"Wҹf�|w�0 ��l���+��v]v��V�Q.al�W�<]g��G�ɇ��7�� hRqw(�$��� ���$'7䩲n��s360��H�?�u���k�30�aW�x$�~C-�8bwʽ�(�a�ފ�1���7�h@V�,�0Z���PpGs��,��Z)22(B]fg|ް2�`���V���ќ��C��t��h���Xb��d�p�� A~���_]�줫��b���`�@g���4l7�of���rD�h;�#���������Hӏ��zu�aY���P���~0;]d����&�~�):��{tA�8��^��oa}Nwd6��,{�s̮
�Ж96>k`{D����S�w�'W�|2�+���Pa]t0�)��ˢh�+3�[@�-���J�@�-(�i\܇�R��5��[P5{b�vLb�dx�����3������6/��֧Y~Ű���o��<�ϸ�s���?�6�����d;�Z�V>l��;��2 �h�Q_�mbF�@y�;�o/	�n/��"��|w���1��N�+� �GN`���9�?�G��uc�N�2��S��W(���`َ���`�q���{٥Y$�I��< ����۳,�6�|q��Z9.�B�y���/ѻ�}��r����,���ᝉ�<� ���aN�oO�E�=N=- 5�)'�ey���<K�(��r⇛=LX�{����^�l���j�V�Wy��Z ���N��^|¼t��Z�tD#ٽ���������En��f!%�O]��$c��H�@�D��I�_t�f��ᆽ�$\Bá��ʀ�It]s��ܼ�z����A�s���	,�sP[z�H�Q�m�g��}u���$�@9a�OxZBv�މ�p�����bBa��J%iE�(i���F�8al���a
1����%�zxw,�7ғ�N�!�F��5u����O,����h�^5��r,'��1�\>/��+S�3�mS揞��"B�#��2�-��י*�,};/��M�h&,ՕW
T�W�f��+,i��X|��Ny�PAy����\Ш�MY���|���X~khl����o.4H�mF'���=�u��Z1���πK�V!LeiX؈yE��!F���p�8�mX���[�W%��Gq:��m�)R�m%tB��>��W�ͻ�,����n�z��%��U�e��SɌ�а�쇥M�h�x�v"ʶ���ڤp��Ao�9??lb���,�|&;�#ް�J|�i=�}�i��	�7?G?Բ)9����X�3WU���1��q5g�d��� &���?t�G��?�֫W
vG�r�DM���<)���|3�, �%�46d*�_-
�p��J��2=�b�} #�� ��2�YGC���y�/N�0Gh^�@��<�4+�<�7�]O����Ϗ��mJ=�WWXCM��1W����fF/$T�"�����S��7x��bZ0��m��%jjN������+K�r��X��Ht�&�,d ��9����g���q<1ȇ�X��pȋ�����J���_>�(Y1���?>C�:M�7����jqiIM��y�������ӧM`�Y*Mt� ��a[ꡚ���]���u��G�>�"���ϐ�RRRX����t�40��5���15eX��KSSS|=�N��i"������n�;3S��8y`ķ���أ�� ���5�4��n5ӹ���_�����ٳg��l�:2������S6=����Z�za��vz|DD|*�:����S�:����K.�@�� ���[�>�������J��ƍPu�:������:������?I�.ZR�`�UG��.�R���~�q/�g�Mx�`N�L ����y�u@ ��@RV?���l�׬��g�bb�	f�v��E�K\э������3VL�:��~����b�VC������!�İ�Ț�z`�4�����z�,��4�!|~�:�����K�����6�x9c�����bN���~:FM�+��kk�D`����[�/2K����M����©{䔎ԅ'�G�q��jWhd��Em��`]C֧i���f�����!XX%�*T]P��ǿ�t�����w��8�^.�Y0r��/|�;<b�o1ٍ��j{����B����sB���j�g�ɮ��n��p
/���t��yPHy��=�ɯ�Ŝ�:}����o�pW�g���l����X��eo �&�����K&I-�ŕ۞[8Z3Ʈ�P��)ϧd$E�!�2!d�0|����M�����1�1?N�h�:u�c��!Ë4�={��'��}j����w�+����ZX<S�k����Hj4�����9�_��O��������8���{<]�H��p1gVhu���M�gB��F��=�-��M	�N���>�4b8�������/�.���7�f��_�`aN�U��i�Z�c5z=�t��!�u�bX�g)�\/�b]���l�\/�#��
�u�2��.?�=@d��u�<�J�����~(o	�]����!jM+�B\wLmR���#���Ko�_b���vcR2��^��P��?����-����]�8�(��%��F�b��'�&�a��ȔY_��Q�QT����qXѷ2���#[j��+�m�U�aK��Iݤ�@XG+�2D�?����"�ǔ6y�P�;>�>�e�q�ћs�#������z��Ϊ
�˘�-��+K����76�0�������5p���Oh)�~����S�AE9""RN|4Y�#����!�Va�LPm#ɍ&���ݱ��!�,�r�x��Ҫ�6�������~v��};6��d`R"�}b�\6��*�a\��O�������\;�����9u=�؃[n;�k�n��_�;849��V�����7�/��]o��γ h��G�cG�c��R�����5�2VK
T���;xMh�ph/q�����xF�,�ak������d�#FЫ5�����Ԟ͘c���qbw�DzZ5�v��k<�������.���\��9&�&@���ϾS�,j��g(�/��q��L`0/QO�&񣍻��S�(Et0(+����ȣ�q&z����~�`;h��̖*+�F����|�掤F�: }��i�x�Ğf��gi�Z9Br�u^S�{~K^�d���":״�-�ՖM�=/z��=����Sox�f�;ƙ��KD�|�&�
���s%f�f�a��h�҉�&_���nrm��?Oh����kg��8E��a���JgS����$���7�5��|�n�ۃF����tN��ċ����Y�p�~�\����1m̔(3��L6*�����_m�E(q�y�6�OT��lc5}\ kM�Sw�J�o��I4�o�#E�� w���w�E֎��w��d� �Eҏ�9�s�c��$F[�G�'�z��ŠE�g��3��9����X��ar\W(�I9���)�/��329���<�5E(FoL��'����Rp����b�nSw��a���Ԛ*q��w���/(,Q  �'��ߵ.�jK�(#.gj���:Sv��N�!{]q0J��w�����u��c���q{�`�e���N��byJ�\(;u��c(W����qE����9:��ތib�J��\�|՟9$tt����|驒��ѥK���ۨ`]�8�S�8�;[�;�g�є��:�(�,����B��T�nl���ұ�}�ٮ�{��J=f������/#��/C�����~c����(G�׽QCw�/�Q�in�Xɨ��h�i��!3��1�G����H��SR�#ם��z��&���&Oc3-?��)����q\�͗�h,��N׀2�4���B�L�����/�Ϫj��C�0���/cK��������\Y*�x��K��HG?>��zzh����ūV�P�b�y���[V��bg�4T	���: "���a��.�J�Z�a9$Rz���.#��<��>=�s�Z�n�i(��/,t��G�����w��r6���OX���f�ע;r$�9B۳x��`3YqԸ�Ui �)���?(;�/���62�.�G�������	Fꚛ��4�L�L�H���yN^�+V���og�d�k =$�h��z���M]U���T,(�&��O�?s!�<�>g��tȚ"2�o��'.�U�aaCL~��[߻�����0�6�q%jʔc}��≧���L
���G �QҜf)��ŷ�Jo�lԌ��i���.:DS�8�җ��\8,,���@'�:܉i��.��$��ѧ�����!*F�Ŗy�j��k�̈��TV�޳���c��+���ruԲ�s�<@1K��J&��>omz��R/����O^]gp[�>�<���e�����ܡ�8^j�ZN�y�xn��c���Ԡg��H�����X��~�qK�I��:U�w,�$,��'m͹����n~�'���\��7��Ὼ x��ɾmk%�S�y?�J�wN�[�z�MZo�;B����K��zA��狠�r���H�ִL����:c�B�7��Ew���*��S�^�wiI-}��HE������[.��x�_�?��j� x�_vM���Ϗ2�c���W�ڛ� p��Rc��������:!yU��Ax���K�Q�����yhP�jj������K`a*�{���
�t)ʺ�����\&��/��u�gqG9�S~� ��1	#�>�;�^����#.�L�F޷�L6�Չ����i`����.��@��6?�!�X1��P��5�{%t#3+3�N�gd��)����墜"�R
CB�W���3l����P�Ӳ��xmyQ~J�-�BǮO�<��s�y9���MK���k��������l���f~��ɇ|/�����˾��\k�1���'�w9�Ȥi)�u�h��%����r[:�G�c��aRt%�6��w��$�ܓ���q4E��5D.��*�8h[޼�� 4 h����ђLʋ������.�+�����[$��&og�PN)ޗ9lq��3��f�a���m���j�k���.!R<�`��g�M��ɼ��L*ng�-_LCX�שc�npL���{/���rc�km���zU����.����M��Dr��IO���:c�,�z8��}�c%[��m}ֵ䏶?��{p����+e<􃳂m�e���V�S'�-�PZ�3�%p���N��y��ژD�"s�ƹ ah���%�z3�~���X��t<J��gU�a������g��O)�ѫ��]�W��QuM8�l�����6���+n���zp3[��25�D�u�V���� <�i.q�m����Tf
h�d�z&�q�������Z�	��M�7��n��ϋF>��'8��[�����~�x�Xau ��/<34���J\nߊ��;����J�7w��ᴿ�à�u�GP���^�2�u�Q9Yّ����7 ���R�gMUy6���lL��Iq� ���Of~d#Sq,��=B��z��aw޼�'4����ڡ09�#�e�2w��u.d�v:�F��Ε.����Vy��0�Á۸{㍯��3d��5�%1��gv*ѳd�B�OA�mN��ǡy�:�Nɽ�%��.�Ƃ��O�˼P����Չ'�_[b&Q�6g�w���m2|yt��d;Y�1���ҁ+��ʠ ��g_��y�}��Qx�p�������9���qV[fɢP����(ܞSRw�W"�9�eE�Po���9'9����V��k`Z�����h��x����A˱}�����D���a�|��I\�����Q���6�>�>]]1|�uN
�k	����ѿ����  *t�!�L�ֽA)��Z�X���uPl�ס����!WV_HI`C���_�$N���������U���݉�4��Gh	ҷj	߇KЀ�p[eX��ߎc�׍�K�Nm�%,��TjBN���� Uee'x_��#?���'�X�Nf����n��>���+6�S�ί� �Ѓ�SlxJ ����-�����?��X��u��B�Dq�R����ӚQ�,��[$���,�,տ'�m (l�v�A�Ӣg���kJm�\�D��d��3�C��f�[�?���a���Z��W��H+�j��7�����f�����$�+�+���s��8��z�)���������9�';l�Q ^���%��4Yi�PY՛�� ǹ,x�;�<].*��1�𳔝��Ű���T�=��F�����̹��W~��u1L��L��J{�8�%9��p	Զ� �T�Ib�,��i�K���.�,���}f#� ��j�f5���ؘ������	�4�Yei2�=���N�_��[V�(Z���b諙Ug7��J��lE2dh�[̈Ғ:uF���	Alt#ot���9�Pq���M�3c��b�G&4~W~�3?D��P7�1?����M���ǯ����9Z�t�J�S�9ӌ�]��' ����� NFZ�!�Â_K�P��:MϨ�2����0Q�XRX�,*,Ļ�ϫv�CK2a�����.����Ȩ:���	��[�~Z�~���Ӵ)uНB��ܼw'W;V�l���N���2�S������T�{y]Y(]���2�r��7{�}�(�3�TK&������ �$ZZFfl�2�O�0[>ۯ�w����FZ��ӋL���4:�����Wz ���U���hr��B�ׅ��N�'+k���0;5�¨��!�e�_�0�&�c�@Э]�_-4�F)~��@��bJū�U��|�L1|��%o��rA��ae�H��k}��gs�9��K�E����{k+��oNC���L�tD �%����8]�:�?���mr��V=hes���%H�N�ܜP�x�`�J-�O :��44}C�7��
Z�f�Ų�H3��fծֽ���HyI[/�ٲ��t޸���>0O{|�6AKYd(���K�@5��j�ң%{�O���](�6.LC�,��z`��R�U�Bsfa[�Q��EeMk�iO���!�$����7����|�A�z��z��ͫ�\��-\�����:Lf�8l�����H.�}ć4480�B�e5�f�ori�z�TA7��ɾ/�f�Z"���j���U�5q�C�P̡o#�u	(e'��ߣM|��m/ޯ$���S�ݠNܞ��Po�r�����TDc���ω\���V2��i����[K��v60�|�M���e<��g�6��գ3n�	]9ȋ�B�譧B���4>Ḋڀ�;Hç>��V�Z<�p{2�xptxГ�`k㫢J��~O��Zd�X�l���GpH�~��6T��
F=_HP�q�ؘ=;#|�Ժ�� X��
�KͶ���H�"��d/S̅L6��¯���Um˚��BS�n9�`���Y��RtPl����yM(�x_"����� ��ǤQ޾���RJ�	�8�zLo������'��&�Ͽ�Okj�p1.���������!���$m�P��kQk�!p�rhY�/���做�Y�E�lV364�3�%�$RM��]9��>���Wl�ayh[L�D|���b@����/#�z^F��.5�D�E�@�^LwC<����~	Ջo�STu����O_�Z�y\��ҭ ����r�d�TPAiOtQa�d,�u����ox8��҅J<;�7���	��BmG7rB�>q�3x'�#?��VW��uS�}S�7�q}�"^�o�����h�j*K͋�7��N>����`��jB:r*�Iގ�t�Xޒ�ox=���W�dT��/E4Y��JK�g����cCIiE�V0V��'`��z٣t� �;Y=��E�{���%326�j��w�&����:A��s�c��B�v.�`/�~.������>3ut��(آ^-�����"{5���O�k�߈ S�SGcq�P�����Õ��-�m{⃱� O,r��}f0/0��a� ۈ�^edn��+/JA���)�q��c=�8v�N��DXSS�DE	�������_)v��z�mo�����4��('�iQ��kz��� ��C���s�LE���r���br0�JuC��\{@���~;S�<����#kkkP��I+Q��vg�&�,���8�U���^Z9ʀ��]<"%��sGz�y�)�p���L�37�㔇j�#��j�"� `f�s��~Nr�}�(�����9υ��ܞA��ɩ� ;�e�P
m��,LQ.�����L���e�k�`=��\��cL�`�>��/O�G�_�:,4�߲��U�A�w�{�J�Nqhct8|϶��e�����긕�W������$.�fI����T77ٌ�=[^���&2d���w7� �,�	T�C@5�w1�:��G73�p����6�<i�w��׵%�6{Sw�T��8RN��Y�Zd��w�i��$������_x�z��t�LZ��B�8�cSSM����4�TJ����R�΂Y�/�� ˮt�5������lU VJI� 3�?�Ҹ`�z�L�v�U1�X�Y.[*���:���Ϊ]=$;z��A(�Qd���>j��V�M\+B�!�q��3��'�����ka̺�<��.�`K��Xg��q���������in��kd6ʹ����"����v���o_��Ӭ�"6e�3w�+綒��$W�0e�bN�;tNh�n
j\�1����oؐ��PR��h���e:5��Ú+�БԞ������ϸ�����A����
4�� ��D~5�>����!`�w�ʕPVڷ�,���L�\��m�m�RK���ճ��fz}][f�\@�JqI!�.(~�$A���)�� �fS��SQ�f-�Ƽ B��bk74���}m���Fn���7۩�4�u�@�V��Ե׬��6�~�*���_�犏Ss�?�,_e
4i�Y��+�2��@-3%~�-l$T},��l8�r��I�^�=BU�:C�u��Smm.�w�瑱�/e��7yҿ�I\�t_�/LZ��p W�,�l�Q{�)�EP�N���x�%�c�����oF�n�[�%/��y+�'�,��p���(3N�l�_?:!{4vښ���i����kB�7�� ��̰�*#�n����@ܺ�0����o�O��bߊ���WĈ-�]�5M�#�6�Z��ݦ��#��'-�Պ�Vz�󣏫��L�\@��Jn�ϡ�Tt�F�wW���W�6 �_y} �[����B�x��� /�wpN}��f�(O@��5��s[ӯ�B��&���}xX�$���T�4#c����Ẽ'(���&0�,F�����1�@l��Q�Ԇ��`9)�Q�Y���57߯珤�Ov�>��Vj��K^��Zl��oV�&�)\�`���"l��ky�ܜ�$C�Ceޙ�^O�Ϯ �.\�).�t�=n' �F��	���s#
P�\s���M�#,6�� �O)·��ty�[���-%E��Iӗ=�����Z��g>��Â�^��8���r=ӆ�>B���,D�����3e�����.��8�V2��d�#s�S�1���u��ΰ�C͋����;�aCc�T� �!��
�M�=$��S��������R�ƋC��W�f���ke]��}��S��yn��5㉌��?%�&�(+���R^"z E������6��3�2�7�
�"����I���|ҕ��8��7�Ys�:s����:1�/���7-<gvO�v�� YD,�t�����W젉�/" �����a[e 5R�]�� ?��
��D���
k-�WG哃)�!_?ݣM.`~�=�e�<L+�Z�9��({�Uy�T/sOÌ�N�T��4���eA�(��x�FX����I�<��qr���/��y�`�j����xpa�A��۫�qX�"JK9:Q�+bذ���.3� ��4�E=��V���v��F�z�K�>��#�0�R�bt|���,!Ҭ+��7�1���.	�S�������C�]��g������FN�-_�1RpU��1��o�k��zg�y6ۇ�ֵ+�c��[���Y��0��rD�xT�Z~�67��A�D(�'�>?�t^}��l�����<����E&�XJ����I{�/#�֣jDr�,ذ׫>\���p:����H�J��-���7�� ����3IM��(����`�̬�J���r���{,��z��xp�����ΞQ9�)�WW�yi��Ƈgp����0��\�G�gb�ڵ�;���W��cۈx5c�~�v�}�lP�������qR�y�w��u������R'�:!�g���QVy�/�~ݬ8|��L]
~ɡ"�,��]����S�K�[�t��\��=�nm��3�F*�i�
\�{��j�A~�F�4D}�����:`�y���1�JA���=��7n��#2|�>��sk�?��N���DX��A>|u����;�F牡e�	wY2_ `���A1Yӟ3�G�/���'N	
�����k��x�MCꔕ��> �>}?q3
��~���h���zy]�d�~������G"�Jg�`b0������--,��;뤾�e8�C~*N<���addds�e�h�_F�g���z��?1�Dm:�  _ 8��ܡ��{��J�R�G&��a��*�=�i�!�^�M�%���3�8�,T���Ւ"�s�<�}qcC[ꬕfc
��J�&��R�G�Ŀn �:CX0�y���l��c߯�K��X�X.�&��"O#2��G�%?��Ӗ�����57O��~�|T���F��7�G�Ё��%�~{^܀����ڨ<���-0kXJ�O5�M��u\m�۬���|%��b���:9d/P��X�p�� k�2� 8?X�M��3��L����&�ik��R�����Wןؓ��<N�3�B7�ϯ��x���<d�Թ \uY
t*��<�"�-�-a/StY��n|Xn�G�d�����+�{}}�7A�y5�x�Y]�|�,m	��>Z���/x�%�䤻O�s	�ܳ��ǍٱXR��V�y���U�����P�A鼦���5�����Q,oN��W����_�<���<�������@���i����g���Wn]��_:OU{�o����ЫH����
�*�.\�iiQR��n��6 � �ݡHw�t�t�Hwljҹ�t����Ͻ��9�Q���ff�����Y3�1<,?�L���b��Y����8_		���y����|�i��V	c�n=������2�$��ݹ���{�;�0�J���u�� G��[�������o�!@ۯX�gm�H%�(>�_=�!�?M ��-a�k��⇴��Q��������,�p��N��������f>ϓ�4E"Z�4Xy��¯�ޞ(������N�{���W�O��7��3��<z��G�ׁ�M%������\�$���[@*��惺�L~&h��V���~��dɀ���ٙ���������z�iN�e |c�q~<���6]gg���ݹ��0k��d�W�v���ᰝu?P���,/��:dI�~��_�`���6��i�����ʊ�u��E����"�ճ1"�y��G%M�'����ɘ�2oY���7�ܞ�9
1��������PP��h����4I-h?��w��ɜ�W��QiW7D�/8������~�T��H��㜳r��ؓi��F��`���k}0�Z5���r.	���, �B5@Ā���1��m<���	F�L��3�j'�������68O��
�"��{�o�W��i�J�TT:���2�ʘ���223�s��D�� �������G��̬��JDXXUUug��墽4;l#eEH��{${
i*��4�Qc�j��2(�}���jf�'�?jns6�`�.o�Eۗ�3ȫ������V�����{�Ez��1�����cBl&�CF4a�� =�,	ͮ(\��e���YG��͡�.�0G��ݭ���r�� �:��]5����o���gb+�;��L���7A�&ݹ��ʿW!}�j�x	2�;:aҐ"��7��'���Wu���T;�-�ȽO�_	�lL%�a,��FW*4#O5�v���le��f3�#`���~W��.�����s���?t�V	��]�`LŻ�+��R� m���O�l�%"X��؛��¦�; ՟�4�p�.�tv�F�p����)�K��W�Ky�c�k���I�������x�bzh�5�g� ~��m����`�?�E~�а�^�\��ՑV|go�l�>A5�<��#�c��i6<��n$��� ���0�mI�f'�=RO> j�;0.#�褙�G�ytAr�-L�]7��,��[C��0}�A�21,��׋̃�R[uͼ,�O�D��9�6�@��o��+}�H��x�({ܜ��U�f1|�W� s��$A����o�Bery�~��(c�*�a&�ru�0H�8��/�;�|Z�G m��<���Gz�,<%�����/*�'���
l.���L���^���̼+w���w��o���?]�Z'��^�9�=��[��ͷ����h?��~��C����H���xϳ���쌘�g���� �H����B��~�ׄ���7�f�7�$��͝�������5#��^zw��D�7����J2���A��b
�]g�����n�ܯB�bJNV��[��{]֤o9�F�{��Z!�"MMb�d�*�KR�˴=5��OB;k��8z�����[�]����t:�o;�%>��σJͅ���-f�����ۑ���̃MT��|�:�D�#P)�����,�3p����������`��	��2��^������v�9/�:�O�6�v�c�mS�|��w'Ap�ٻ[���f��1������7�RbC4D��5u�Y��~Dϙ�����A�����yʲb�q}
�? Odf���Zq3�>]���݅���{-T�
/=��x���xWo��>�	|�f�Ҩ�9���J�����0:psi_y?����e]�5U����%��]򖋇��ޅ^��e;U�k����:�� ni1Th?������I	
�Z�0�B��d�X�Qx�W�<�:u"��zJ<0�f^�k)nu	"�r���Ei,���_�&A��B�l&p��)���'��/�^����:���.��e�j:���ϳ���vTm���,�:w�Dޕ���qy%�.�����m���D�:�2Y��ƅK���<oy���4�ʮ_�ԛ��HIU=r���ʌ'���Ϳ�����L��x�#�x�i7	�S���&�˖�?�I��C%���{��gG��B�DTlb>VE����?�ə�t��Y�<�����,��==�}��wwT�BF��h�?�S~~��8F���O?}Ԟ�3h�[�5���/3�o�O�Hۈuv�Uon�s�������B�(���Ud�'��Sl�#�E����J��C���P��?���{7rjZ���\o�Ѥ����lh`k�,6a��"�c�k��h���&�o�����]U�W!6Dō��\}\s]�.E� �p�g��x���bn`��S�;��_������!?�Z+y����pv��t�<���٫B�\�+��Qׅ����D�;IU�MV�WOX�m�;��?w>���Ru�0�����,*�;2��~��ŦB�8Ϡ^���I�>γ{{ԣ��9��a=`8U^�d����������6[?p�X�f�dQ��%PeG>E���{2�z亢v�y徲�����j?[��4�y�A��h[Θ,+͈c����ԏ�Wl�.�������X�)d��K���a?��Ro5�"��A\��?j���\\HLn���l~ߧ�Y]����w���射شVV�%e��_W��_���Y�okwTR���=O��־ۼ���������>����Ɣ��ۦ�O�P�$��Z��j�\~NxH�6c�v��B?�W��@�!����yxe�����i��?��b�di&������p��4�q.�)��^��ﬠsAye���-�o������Ud޵�Zہ���	��)��*&4��H����`�eF$þr5{p~wY~�-��+�M�.����r�?	��������\�s[BR������؟.�P^�|�3W���� �E�}��r�����~+�����*'���ҒO��m_�?��N�nԦ�sA�c֦��W@BJ���c�7�t]cs�VI�w���C�Gū�24��U�H%��>~^&���u��,���}�(���\�������Ib��# �-�7��c�z���+�|�Pez��J��H��������� ^�F������?���
�s+���}ί>㏁7�G���J��d���D�g�&*�J�9Ѣ8��c�t=��xK���3:`�&0̴�������L:�_��r�*�.���nT�<�!���n�s��1`Se�����J�SK�R4�?z�"�ǅI����b�<y�9g�`Ҭ���&� x�E,fc��\���ޤ'���f��B&�h$�ҵP����4�#�bY�#�9���&w#FYJF<�cLLL�vI��m��K�=���#\�s�[;��ô[M12��\�����E�.�f�Sֿ@���m'f|Gܜ�c�Ȭ�lD�ᄛ�Iz�>w�C��SK��6��r2z�ޡl��VVRd!�\@���D!�����b�.�	�h6 qLG2D�9xzk�]�Mz���_�C f�ɕ�&�/�'���LMMov�Rds�R� vqs�RZ]��M�Zdx�d�>����`�|}����Q¿l �yJ.�0������ؑ�˃^m��=�^�ӥ&L�z�æ�f��u�d��bI�j�YcD�h�u|�X�{�|G�B�tt�<�3\7g����î�ꮭ��5�PPX(����o�GB�Nj����H�߰�Q�g
��;@�,Z�hB�fL��b�Re"��g��x�%\�;��!�H��{{t]g?�����+�~Um�T2go[�d6V�@o� ��d���9B,�y��i��t67�����'"N~��������>��+�ćJ}W�M�u�D庛<�����h;�|�A?~)��ߘ��Q��:���2���<�ӷ$��GTt��c�\7�)��$�R1(�@�P��ED|�:ْr��D�M�*|32(��`M��̃�&$*{�A����O���_���#n�����`d:�v�7_K\e� �����=�'��\Ć�Hg�Ҙ�?����qq���5�ۂ�L0�C�K�e�kͼ7C�v��q11��0v�c���?8O��0X�ЉY��f����O��c����i�B�I˳3A��4�ɵ��9?�+�Ǿ�\�͓&)l�<	qA�C��Z�l����j�z���{c ²���\}�WOǗ�k,�+�n��vg?�X�
 |Bge���_(�ԛs�{�er���Vh1XH[v	h����,@��\�$گث��QTV�F%wX�P��)&X����P�)1��Ff���iH߱s���R���O�U�&�YD�f>�)fc��l���b�����r��{H\�0!��ͨF���\Gui��r�����еD�@��B��U�R�lR���q��"v���Ւҟ!d�O�T�����C��^�r��{�6\E����M�.u 	��� ��zY9&��X��ǧB�g�����=�IIU֋�H���9�14k�-kxJ&I������q�͍b��x���a�>�����Pm�]����ށ��7�n����P��S��=/O,ۻ��Uڅ���U��ed�\�RVP���+���Vm�|n8mޙ&��ԑ�Q~R����M��B3��_f�<e�^{׮�a���_(d�DK"cM���Kz��}'��l�\�M���p)��j����tYf-9"_��L�z]��B��j�CǪ&�_u�9�q���y^By�,ߕ���VZ���$��g?��џrW�O��{zF��_�2�8��7��[�����5d��=չ��'��PJ�͞���.i�w����EMD��	���/��EE�;�g�i���'�*���}<]�j���� �͘&1������x���=}��i�+{�F�\��1��L:5p|��k�}JZ�>��}w��������k՘�r�9!K�w�4���C\�Z�l�/��3��m�!��+*¬hmm�K1�������\�?�X�/��Q��~	G���r!�'	$���`���?�v���WD1��g�o2����U�|F��@��Vo��S����TS��Dn� w>��T�!��ra��?J�V�,F��X�iS�;�6c`-��H4�H܂��q�`b-E��_��J�Ia?������K:df��L~_J�.v0��>�H�� 2��%9��Jv�Im~>1�z�z̻����N%9�l����b��T�������u��9�!@�7��Pe�c����-�{u�p��=z�z	�^�L�]�ۍQ�x}h�Q�~m�]yN��-&v<<<�J�'�'6�/_J�,x6 �	�"��������.��G�?�`�!�L�����#
V%P��:���N��]&`�74��7!Uh�ȄVue��ȣgc�'��̎��E�l��T�������.�K�d�<H��4�k�Ӊ���C����D�4mֆ��b�;�{�z$q�E���`FQG�W�P14���vܚ�?�ǟ��"�Am0_�.1�v�@���^J��e .2C侥~?���l����)��6Zi�����5Y�`(�6������Z��i{h����w�j���`y�����y���a: R+�ٗp먙o��;W�k��褆K�[F��5����������L����O����3�������rr�d��:1C�����9��b �I�6�oT#в���~����.�\����w�5T�-K�ģlR���P�ЩƂ�6ά_��$��[	3qfy��d?K?	�����-ֻ������gQ�1y�&˦c�i�e'Z����f��>%��i+#赢U�V��_�T��Ts�S^�0e
v����Rf� �6�o�/��L�������'azk��ܖ�<�"�	���O��1�[ؙ�p�6�K ՗��I�#� ����i��Ԩڭ�O��z�~�~D&�L���Xj]�m��5�VY,�W'c��P�;;LEk�8�G,.g*l�6����4hYA�gh��)�M��EԑkȜ�4�!6"i0���^��}�6����R�[U�1����,L �x��c|�J,�
�������edl,�|{y�A���M���X��~���:M'z�V���6�=�mwf)�,~)�]溧mUUr����=b����H@�CN�ό;j��	�gP��*Z?vu�� � S��5Cc�"���@R�U�����[10���X|�	�R �'
x5�`���D{p�~��������Jܻ� ���������XO[��C(Z�ﾁ�H��a�)Wy���Ӌ�!Zh���{ۛ7����wn����xnJ�Qұ����=��8��9��f6�x<y�W6W��k��D �6��6s�,%������2��_>_J|��:�@�	�(��I�V��}�K�"�z8��K�%[� ��Y+��:��;a��ԙ�<�
�3��9��:�[��kL����uvU��e����v��(��)���,�X6�8�maR��ׯ%��Z���>_��q=��4c)"�I�ߍ{J�Bh�ˏ*�&���աI��#�;���/�l)�4�f�q���a�`>�T���s�f�G���q:<2�X�x�V��#�f�X{:�v�/p�Vy���� �Pb���wJ��Z�� ���&X��������;�_t|҄�q�g��:���'[X��$i'�
N��~��:�N��i�'����bmO���)�ܬ+,j%U3;���Y��g7�6��ҭ�z�uבR�?�^}ͬ��خ��Tc��q��.��ָ�Z]_߾��Ml��S���� J�=����B�n���*������|&�N}$�-�=���ż5j3v�pzJd�++Y!�<�r/�ED8gyO�E8s���ԗ����]�eU�O��6�>w0.���ƭI{ �'�����w�[����~��M--�-<L`M��n�� ��<�C����a�(.;�9�jk�u�U����c�`�z�K|�iD茀�Ӎ��k��wu��I��S����0ԥd��i)�����q�$dt�o�0�b�;}��+'R�M���%@�.�YY��3ɹ;��DZ���j�$�4��n�H�y�<>H��ZN)�s��&���4@8;)m{�bp�YG_�X�#U#2T:��*'jfn`_�9TRaH�9O.=��S�虒jb,�ͤ�'�`�,��'~Y;�m a���o�<)�6���TΚ�[��5:��Җ�a7S�K"""�<�<���ɹ�_i<B���Om�.T�.(,Q��Z�@߷��>$��^Li�s%I-ʅ[eHs5���Fۨ:�y`�&�*q�jWp=�T>ބ(�۠��6A�)�i�a^�F,g���Y�������}좊��m|����\u'NQ��Z̖W#�nRn3��Z%�AQBBBq�е�~�ǣ*Sp販'j�lR:�3��j^-�'cl���ۥ-�t�)'��[�U�F9']�^E���oo�'����w�����
����(3���U�aw����<�X�&�N���z�r��=�0U�1I�u�2Y�r��$�;��aqf�W[(��L��s���U�ˮ�ު�X�Z�?є�/l�;��kV\b"��Xb�J�Q-T-��u���$���Sb5��U��V�Uz^��ݜ-�i�������ŏ�31RRR��%��Q�Ԋ8����g��jGEyE�����;Tŀ�Ȗ���t�ȿ������Ww����Xu�'�(�y<y�0������p˺�G��=�Ec �M�'�W%��+��s�Q&+'�Q���%r�j��m!��3,m�Y�j�;~��=�AI�(���"4�쏸[ �c0X�J���l	�0[7��kO-��ץ �����7�#�@t�w����ڴT�YN^�:�J�t\Ϥ��՟-L>��-����X�4U{c:gJ�_?���тMq�y1�����Ɖ��e����������O��6�blIy�v8	i~D�y�դ�|��ж�a��WCJg�׿
qU� ](�/:��}��o�¥oP��f�����bp�HP${����<����N3�1x��j�˛Ǌk��ܗ�g���fK���2>�� �Z(�M���3��n-����Č�j����`ʁ��|K�|[�j��P�n�Hu	��$ƺ&1�#�z<�xf(��#!���'y�S�w��5�#q}+��_p'8pG-��2�l̎UJ�?7��r�[�^���Ț�3��l�#
5)� ��jC%Ϛ�l:�}ijj:겞b�{���ǉA�[�s���RUEŌ��z)�� !n�+ϖ�MG�Sߟ#9F��J;D(����.��.LU
����q���6y�f(��UJ�7�܈QV����~�b�)�+��捰�Z���#�ْ�g��?Ύۺ|�W[�	uy:�=�~[��l�Y��\���ư�&)q�p����g�M� 8�������)��X{�ms��o�e0�8c�r�E�a�H�����(,mV�?�>�HH��3�Vh�͇֗@Zk����E��S/"q���T�����kW�қr��cAQ@�ޞ㧰�}nv ��J����!m������Db�[��|�<�|:4�L��������h��wn[�%*Ė���Փ:�uS �$�q|�?h9��]zh�N��S�G%�+C�%3�)����>?���	�+"=�J�.m�q��y�F�a�k��;�����^?�{��<d��4�x'���}5[�{++|��X�8���}n�#>I�k3�"�4��  "G�nwA����9Q��{�+O��pJ�u��(�2��6�L���o�u�N����y889m�,�g"deh�?�����z|=������Q�qY�0�6J��J$@�aY��߆� �f��)��:��X<)읨2R�R��`�#���§����̓�����vֹ7����<�s;�d�\�p�!�O���pR���tOC��� F*�\�)���fc\ϯ=�cL�*�eA=!�/E˫��v�T����B%*M����Õ��IpiG̿�p�jٸ/:}s~*D�8p��q6�f��/J��e�3K\G�R\�VH��C�^�=�^�pm(vt~p�ۮ�E�gK�X�\ߤ�ء2s��W/Z�,���s�4'K�I(>TC�6�0�������9�6�Q�&��-���{t��F��7�|�_�?����[�z�n������̃��);��n{��������xM���VC���/�����a���=�����Out���AH��u	0(x�H�PM�pN����us��[������"`׃��|��q'���k����q���^��P(��Lk75���ݫx~O����~��ϳ[��U%1�3�9n��2�T��W�+k��wq/}$Q��]�H���h�DN������fv��	D��vhppb�c��^zOOǂ�Ҥ�WS�h͔p'B�e�ޗ���N)��aX�>G��e����k'><�Kj�����|?�U������e�-E��_��5�,�
+h���zs�_�T���a����Y��R�X�|�W	��W�o%���Y��xH~�K��n6oS�r;qx�c��ٰ11}�1t��P��XHH�5s4��uL�\�,�T��O�t�i��]��\��5�e�^m��6��ko�G�A|��.��tx�{{�N��p�>¹����\�NxX9u8��C�m�=��O-�v�"�<�<Ŷ<E���*,�B
���)����sDJa @�9�,��~1���l��|��+Vmr3͖�� 9qr�4q��tg�Þ�^h���X�����d����M9��A.1H�E�eU�����������*�׈A�u�B�Q3�H$�-�p0e��s� _�{�zo�]�}������uXU�k���V���ƭ{�H��Fr��MEbF�Y�����[d:w$���)��PB�!ő�����+o��WUʬ B�Y����8PUYO��ky5Ng�?i��8�����~��f�����������2�L�6�fffX�v5110�ݙ�Twp�kgY񀛭�)eZ���#%*���h��h	)Y��=wݦ�򦩳8-M���a���-�\�s��-��Ln+�BU��m9yz�(�]B��m��ֱ[͛�\��Ȍ}~�N�z����d.��K?B��K��&E��͐ok�a�
�6#�[Kr3�@�{��/?����6A�ynu��<�0�f䃒��v��r�9�ŧ���UM�������z1���,mT�O��#s�J�4�����V˶�j6�ѕ@����q��7<�����f�K�2%C_��밪ss��1���)֒�At�\�>7��@�e0��C7	�U�Y&��Y*H�/9B���B�v�	�-f�4,�:v%V��{����0��8;p~��C�*�T�]�i��@���g�+[~f+������`&ʅN��j�F�*���*���M��[&�����͋IBǔ�p�-Ug"S������w������d�̰K<P�6���E���,}Z�)� ���H�=9�[�ti�(�S��iy�U!�W3s���^L�:Lou��u	�H�T�vT�R�n�9-
h��ʇ�����pFH��~CܢPx�b����)+ҙ�H�ѡ�Q��H���*u�zSXi'7� I2��������3Q�\�,
i��X$�Y�Y�� ��1�Y$˹��B���Hդv�ӂ��-�:"wSs�L<8WTS���&�b/�0'P��/���%i�p$��| o�صXC���@Nq�#�%��J���R|p���3m/��4���e���<F�ߺ~>��U�"m^��+�E9BWg�?�N
���Y�֠���ܕf��}D��G�-g��|iX��8�bL E6A��FN_�m�J�� �{��4?�+��.��s����`!djB91+[h�*|NthߚE��3�P��fK`�h�X����]@�ި�z�O
L��yT��[B�K��&����WU��y��s��������2[��(JNT�N�;�g�ș�A'�rgV�.���ͼN�L�vؔ�G�ݬ���j�k ����)��-X�f-E=a�8����R���]���������\S�@ߢ�#�����<A:���Z[�>�ZI�/�+�u�T���>�OZ���<�r�$����v����3�h��:�+{W�S���	�bS	���r ��I���Ղ��.��첕�k?�w�:�>;��������Iܑ<��S�s���4r8��������|���x1��F��}�Di��L�W���#L���R���4ΰrX%��@*�<Nq,Lv�`�"�7`��Y�_[ѫօ��]نϗ�TRGi��;��o6��H���Y�!r�fMq��k�
�{�U�`�fA�!F��)l.�kaS�":�y�v��m.�||�2���0���-s�� �/�Fߐ�o�-T)Y"�[6ww�y�i6��\&rX�R>I�}֌	��M�>�h�ۀq���d��%���N�˞��ރ����֪�q`R��+E�.	D��q�@F� $�A{�D���q������i��-t�ZU����PPF��E���!o+2)0�-r�R(j6-�ۗ�>n��|���D3��À3:@S�Bq�2\rU�!m�] :55��������EW���ЬL0�E|��v���?6e�*�{������
�9g����=z+�S2%�\t9P�!�:���ou8K&QG��&[*E��:k@*�m�R-�d�f���4�hyt�]����D�TP��z���"y3�b���8�&smmn2󠏾GT_y��A�o��*��@؜�:��x���*�U���:/\sϗR�Oh=�P���mSs��$�tD1��G&����ZY�����_%H�*�B��h)����rC�^[��Ig��ӓx/f�=�XC��$�$(�*r<�pU�����e�QF��KF��W��e���@�����> S�]$tJc��d?2�u��u���|�\$�z�~RP�}/�Vs���
DC�J'�^׋kT����8AN��40�h6�ظ�Q��Zߓ��.�O���<�e���]�	��(�s��@�n\��kaGg<l����f'�u���r�D���b-I���Rf�C�7p"y��n'�~������Q��0�C����a�e��{?�k�4�g��ە��hn:�
�����{��.JA�dp��
�==8O��!ycc�U�/�Ү��q ���2Q|��U��7#�z���R�bql*	w����)�ө�߭���w�������^��?OTY�Rw��;mr��@����}�/5('�V�m�XF� ��l_��{J(6�H�;���Aj ��rRx���>gAM3�0&@Q�!?�D}>& �����s8z�r\f�xc
i�������?� ���<����&���!z��~ޗ�(�!�����~ǂ(K��{	|�����z8#����?0��1���8�]) �;>��(����a�I�@p�w��ưK�<�7C��f�� ���B�L���R8��UؕMܼ�y��!=�W6ujh��[��O��O0܀DUP�
}
!�,�Vm�Q2H�6���-�h�J+H����i6�?"�v���I�_k�J;�ڮ;t�jf�1>2!�c2|��J�y��K��Ιf��Y��)2�ҶA�!��F�*/��s��+A˂��'M���l���~�@�w��<H���qg��v�����F���T�w�#��Nn�x62���gO�׵����BU��Ft�v�m�����H�N�7��'qh�9�Ĭ��������r8��ZQl�u��E���8���0b���|kf��:/5�lđ?�X�(hЙ+y������`���:��|�1�:���א�`0t
D�տd�ʨr�!�D@J�^x�+,h�1�\Dev�W�'2:r��A��ߖ���N��94:88��[��b�Aߣ��x��x�X��ƣE28lE��
����\�]�AF��?��9��.U%�q/��@B�_݉���1�2/`|6�Ȃ�����]az����|	�N���	�W���{zy�N~#�=Y
oO��6��F��Nғg�M[O?���k@Y���ЬC������������|��qV/��4�P��#��(HY']>,^�.�GwkW��yq�#_�Z�GZo�_�\1��%�>_^�Ϧbh�R`^����ܚü&"��?��x*<��c�����vi��#�/����0�LVb�Y1ɚ ]eNNu��K�l
 R����
�Ո�����G�b�/Qa[�z�z�k�]C
g�*k��t�qga��X|��v�]H��" +g�u�����ɱ^2B�s"s��/n�P��m�!��3M�'	�d1��{�q�}�%����P���ԭ{��9�y�d�\Xyꛢ����`0=5'(ٌ�� +0�o��^(�b�Ht-B�o�<R�"K\�L��h�ɀ�|�HM�/�tߪK&��!������i^7.s.�)9ŏ�Q}c��4߬w���F<y�VV�k��O�$��˥���f�D�� �	�
��vX�F����[ϰ�qCDʂ-�J�;/c�Y�c�fJh���Iqw����m$��
*���
F�Y�����b�$�h���&QÇ�N��N�界'�;lIj��0�ӗ$X/_�t9��C��0T� D0f����)���C�f�F�*�{?ࠟ�S[ac����ԯ��2^����Z<÷�-��7��(�~͏�fz��!�A�s�+������p�Q�H#ݟ��Ujk*�Bkm�ry~��U��a���IV	���ң`�ܽ����2a#��V�}� ��~s1���W<5�[��,�@�C%��J���n��#vm�g��8t[�&��n�m�H��H r=�OuG�!1E��Ub�+���1+�l�m�	dp.]�9�-◒�{�M3�i�	�ǻv@�_�w��?�K�5>s�~�<��"�F*Ho;S���<���G���Ur��=�V�N��dK9���O�OC?�0������:�>��<�R���2|5I�����l�����#ۤ��ފ&�˕��x�M�����[���X+"Ф`����Ԁ����}g���0�#�����
<�>��k�k�ʍa�zH�9��I�����OQ��2)��
&��i���3�	,��?�a�� k�Y�C��B��$���d�-pRʓ���.�E��3� ���O��� ��a2:�M�z7e��Ca,�Oo	���d�l�B0�����-��j�.���nT�>i8��VEt=���<���P�I}z�I�_��/.��N�.��u��x�ÔaLR��D=��-��W��pRӱ��e��(;��+��	�`[��� \XB�;����Q��+q�ۿ�q|՟y�W��͆d�&T{5�P"�[)W�;.����&��ʅ�RXFL_�ig�?��@H���[1o�#�������?8���`��GD5�[��ζ��v��6����X-Og^61* E���4)�7��:�]"��_���<�ev]gUJ����U�r@���p��+&H�IB�e����"�O�#��?v�P	���h�O�W#)t*�n���<x��B˕6�؁�>NiW���'w������v	�|�7���"R�~nxd����9���~���)Hh�"?Z�n*��*3�N�j(vb���ټ��t����{�.��F���i�`��HF��|-�b�.��J_6�Az�q�E���ZMڞ.#�Y�vD@��E�_2h�M���?dl��A�Lg{���C����B��-�h����>R8����r]���2/�+H_d{F�n$���@z���a5���0�������X}��̉�5�cp��m���ÿ�[��@��)ֶ�Y�)�G4�{mk
�ޛm�Dh,��Ij�

�JG}�/Q!>��o�����|����!�D4�2����v��|�8s�K�'�C@�O�E�i��@<� dQ1'v!x�$�RknZ�0NS�)�:=T	|͍�`b������}Ľ���ZzI���)Z�F��w�IrXd�]�Z�C��q���A,�cG<��!��{ܣ�*T.����%W	bͦԨ �et �B���r��-�j}�:��c]	높�@·F�o��Q"�d�����{�?��;(���1Tك<N's%G�g�1�#��l���ޣ��^��r���TY�h�/<���KI��2����L5ͷ�����@4,H;Ș�)��z�-Qh���zU�8Z�M�_=u�E��T~�faY1���V��uj�J�[qg��1�@�P�E��9�]Ƞ_|~G��*�v:�X-��Ǚ�P�R�����N�`�˗��,a�'	�\�6q1��|ɸ���C�R������"@�[���K�W������W�GL�f�Kq��O/�~ ��|��U���j��R�?�F�5?��0D&K>}��{g#��������#��@�� ~���LY����(�n�X�N��Ց��c>8�pHJ����dQ8[���e�b�~��0��qe��0f��y#}$��:r�}b�4H`28=<z�_?"�y�����t� s���ӓxq�p�+����&HiR��p�������c��ܛ����s/�l}�����f�Ar��ɼk=�Z��h�V�Ն
֦���0������.Yx�IN7������?�!�c�� ��A�)�-Wgs�\#@ �������������ݸ�@��NC��e ?���w�:�����"����"�sֻ�s�!ƙ����Z�x��<�{5%#�5Df�6�-6��ɾnW)m�޽/Ho=]x�
�҃
ec@$�f�xy<��, �g���p���8�W����<\C�p��L��#�qz�zJ�[�0�U�u�)c���뿃�u���7g���I�6�O Ja�?g*�A�& ܦ�����g�T�z/؄3KА�_F#~w�S�ҥ�����=;�_}��N~o�t1iyx4Q�&;b�|��i."H1V4������pʹ��P@��lQ��ޜ�gM�t޻z荧l���\��ԡ�I"݄U:����1���Ä�GHt�R�7�ܜ�9�n�`��˼�^FQ�kd!b��=K#KxR����?��<Щq��,��d��fPi?�7`�x?�%�NM%�b<:F�-���]F�8��T�yO9$���z��&���n�&�D��v���e}KO���F*��=�2��k4�(4M:��5��Dz��������Hi��.��`��<2b�������6	;����M��YI��r�z�p\���v���/:��nJ+�H�������HV�w"F���[cj�)p[��#*M>y�X�4�����%s�d�	]8b,��{��-��}}Nh�\��������Mƙp�����-���ň>�����·�Q�.��-��E�]cn�'8�"�#�ߧb߳��_Igcb�2��b�E�P/ffE�11ύ����������晩V�\*eæ8W@@0���q"����<ٰ2b�(�!U8� KƩN�Fy����bA�)��n|��ǰf�t�8�g���3�5���
����0�����m{-5T�Glrv�>�&��_��aVT�XH�h�b�Q��N�����Yܹ��b��c�A��@������3O��(T�
+������C�M.�(�2o�T�֎%\����#�k�݋cg�6��;�]�m��:�7�/b,A^��v�˘o��#�{~�lJ�hsN����!T�5[稳�wd^^X?�r�.��E s �rw&�cL�6��	�y��K�		y�����E;1�k��L�cL��gO������^��zQRZRQ�Tr�P�_�Qrtӗ�v�@��6n[�=1ꇒ���n�'�(4�� g�me�n�BMBއ��Ԏ�NB[_��_٤�_�jt��a9���{w��E^������k���-&��N}*�B�l�R��C���pG�_pc#	*���(ǐ�=d <�T+#�s��5Ӯ ���#2�!�������.$�}:N}﮶���~R&�ؗ�x��)�SQ����A\�,�W��z|&���l�4��5�� 2b�F�ܞ,����pOY���֖8c^ӧ�ɓѹdB��ʻ��1�7J��C[I�q|�֘�gc-\cI7��e�|�eY��R�`�����u�ch{|�*?��V�؍�<���E�骃��9�>�mys���F^�S`�=R�t�p.>@B���,�<ڃ�����9?$x�#��0{ٕ�?���ςB�4����LF֦��ѭ�TG�d��ۓ>����w���F�q3��kJ.�e$&v�N+͞���������١�f��Q23��l������D� �A�*(�Nif�o�o��eʣcl�HO&�o�zbI���H"''���j~�vp!���J���*_���W�x��ɓ�,Ջr�������Q��M$�;�Z��ʼ�"&vw�ƈdl�68������A����~ɬ_^�zZ�@�{�CO:(H�coe���.��ª(
(*�te���(�5t�(H7HRҡ(�� 1 ��H�P�yfpw����w}\�׺��<'���9�9Z>����ط'P�hO�{aV��"�ы8�},B��ٓ�B>{*]㊔C"YЪX &�-7"��T�y���Em��1p�N�㞜+~(F�*w##4yڕ� 鵲K&�����S�+ccoq��z_3�/w��<c�-�U���=HUQa��2t��� �א�S��/���o|�8j&G������2��>	{9�,??�P)1��N^&�?�8C��
=�l(iQ��������斍����VV�c%�{No��N��iky�<���� qs7k-*'�ɫf�A>�Q�[���'۠��-�»x8��&ڔ$S$a�\/���Ttx��ۃοǵL���-���*�lܙ���nuZ7�=�uzX��⣚��S���T��|�2j����fo�������-p4uߘw k�/�������E|��j0�s���'ߓ��y,V�6���\o��7���֛^�!7o�{�*_���kr�w쏫�A�G7w�����o~��vn޼��cF�Հ[C����W#�'�?�¶i/�@ޞ@��1P�2��ҧ��./���sY���[������J��?����9*�Nr�Tk	�f�)Jct�������'J �~D�,��g�/�c�f�L����.���s���BM1KΓ�:/p���x�)^� ^b{�ɠ��lT>$�pP�M{�y��Oѽ������ـ��o���$�� ��ވ�Å� lP�z8���&�Q3����H��*$�r�3�&6��5/9lO���Q���{�%tU�h�Y"C ���U�6�\M�����i�t���@V���߽�N�W��S{Mpy1
N��/�钒�v�גb�F���Y�_��_0��/��V��.��ʨ/��y����D���v���k�p;�X^Lm��X8R�����A[��-���TrJ;l����Fי��
��Ӓ	�+F�5��s�]��0Y߿��}�I>ȷ#�O��u�힄�¿X����	��~��M/C����M�ʇ5�ɍ��|�*�r��]�4%?_�E_��[2�p��3��v��89hk���Oá� ��ʶ��$^�E�*;G�8I����2 5{��y"V���a�Q�fn{fw��y%�������G��B�`�2LG/��������ך���e�Z�v����X�J�xO&]���FNשP�fJ��3�������%���qÌz�:,����[]M_�r�6��X��B��ĳ!�н(#��"�yV�d@2Y �񩎳ʥ΂g����&�&$ǭ�z���B�����M
�1�"�� _�e�k6������ߎ���z�^�7
�T�ۓ�o;p�x/a20y�v?3�_�l����͜���6^���{���@��f½>��"�?��ގ�(?��|�/����l�u��f�L$��b�ŵ���$����q���06e%�ld� �����������}�4[��N���S��ЫMg}�ɾW��n�]��/)�M!9�oL�f{�AE��l�z02�݁#���8�����O�H c+� ᑺ`m:B�\�e�F?� Mu�$�]�ɣ���T�9j�y�'3�2ǥZY"��i�k`S�
���� ��6Mx^{~N O�(cp�%r9�Y� �Uź�*:%[������ſ&���ń>������Իwn�^ݰF��CǱY�t;'�!s5�5���
�*��]�ܓl�/�#+���r|]'q<tJX�� ~��J�2��Ւ���|[�F�a�q@E�Β�wc�9���|�����@}Xν�s>Z��3�=)��k ���ƶ^�n0rr:}&��)�� �h��/�*0��?F�ɼ��z'Ɠ�F��nll�׽���E�6n��d;?G&�h��a�Ò��"��2�ۍ��(IsVJ�~�S���_e�*w�|Ww|�v����ER4=��҂��rE�~���ّ��]v�a�|��I�4^;��F����.�V�Xu_�̯�z��^��i�Ͱ�u�ō���J4 vjּ��]7�f�>\33H�ϊ�p�D�t��vh�43�Ȱ�@g>*��`u��L����뗁�Uq�	I��j��܁W���lͳe�,�(�2�0&��g�u�+g�� �~�|����&����A��0R�5��&_��\��JX.�*u)e�Y㦶k12�b�Ŕ����Hl�\֘8f�q�^7TY��@J9I[�k�hfd<[S�5��!]��`I���mTT����Iy��?���S�8*���9-3��!���X��^�f�1=
xr��oI��/{Uˤy�W��C�+�/������w����G�Ye6�2C�a�r�]yCQϷA��l'�$ϼT�Ҿ�\_T�닕X�S��հE��J$������ih�_��	��;��۷���o�{���d�UUq����6��wLw$���srN�O9]�h�>�6��c%�-��ځ�"��H&��&�9_0�crWt��Y)u���� ��2�ÏVL��,�hPX��Sl�W��̄���p���=C�7��_��1�nZVq���Ӱ�ͯ/��/����`0Y�V�.�`�j�d����Nb| �D��]0����@�\�;�I�����W��iғ�i&����u�/��G��:)�� \��Z���o<��d}WG��ܝ����Jy4N�����1A�/u%�7|��>��"���Ɵ�)p��prn���+�i\���X��w���rT�<x1�|��-���jW������9�;�gg����?��E�_�t�g!��D�f��|N������SM��&>�Q<����TmS��9��Y��ۣ=�1��R�,R�Jf(�A��C��bh@-���v'��{��n���:�M�H�0�s��'?��g4�mu�hi|�����F��{����v���n�l�	}����ۆ�2`҃���&�
C�Lb���6Dqs|=�_g�Ϫ,�wn�I+ʐ:��v��OM�o�UO��k2�&��s�?�{����d�J&�&�k��ܛh�禨N4��̎�Dr2p����mp�V�������B�t��&�wM���=1�I�E�8��כ�t[����� �<D�)c�Ppڙ>���0�� ,+8�]���/Ee�ѕ�(��H)�g!�9�e� �q� Ɏ��B�r}�ǅ��%����t��!Tj�z��BT����R	���O5b:~ֻ!��C�����;��^���:m~�K�\�3���-��Ϗ*����j.��I�X+(����8u�� ��r����dg:s�|ɛU=ޭik[��zQ��3 ����\��|cϪ�����Y��u�	aO�����BzgYIq�B�q�ݘ�T�~=��]xUM�\A��&�3�!���A��*��.6J�fS~�OU���&p?��?��`���6��J!��ԸV��k��+���ʻ庬�oT��٧�P��{C�+�c<���W[�����gP�-���/� ��FG�����2g%M�A���rKĞ�84;��0��~v��er��� �,����rMb 7��ȭ3�L�9�MZ��1-�`��
[B>ǃt�JH�.��b,*�˸X���%�2���/��������Ny�8�|v����y��əaY�l "sN��(�� � 9�������	�8�-<���,oB���Թ����l&ϖ�^:���ё����(ȎMw��w1y )�]�ۤ0���vO�v�B���q�*`��sS�b�mmѝ_(�~N��x}4�+	��?�]P}����2 4��T�ТU�����.s�K���C�ځ��񪂣ʴ��a��pQJ݋r��ni�gk�Fgg��L�ͣ�Z�Dy#�������Z���s�ˎ���(�����ݓ-<�a6 �A�c�w�FwO��Y�*�����v��E}+�V8�����e�2Gii4 e�����F�ltG�A�ri����H���8oC���-2N���#��ґ�Υ#Q��X"M�kjp��nvE9�k��o�F-������8�U�����!��T�"-����)�c�R���v�uȧ<��
�s��{�
�9u%%�sWzt�9Y˸�M<�(k�6�i�l�(���Ȑ�����L�SZ�o��X~��D�"�a���8X�ʺ�7�~���������/n�H{�"�ſ�N���9/ؚO
۪�Y�\*c�;�OO��� �Mh��y\���߽i8�pz�l'�>��'�H0mҕ�_s�:��t�0IOb������;ɉ�eRoj�㣏-�ǆ���K+$�n?����+�d���^��%_a��*���h-#��E���ץvG���O�@�a�H�=t���8�]Ü�L�g�AQ"`��RJ��Ʊ���d����&��B�/����O�����qո7,���D���S�A���w��Tsv����s�r�����]���N��*p8;3�����x�ˣ��I�uR�\ҘN���3�^�6q�o�k�ſT=Q��_��?aP\����[
����F@�Qu��8G̎!!Ɋ�׬�bd�+U���j~4с	Wc�|i;��Y��S�~<d�K�� QZ����"���0�̔Cw��4�����SY��*��2��s-B�=��o���BM�zj\���lUA�_7�R�W�NQ��An���m��c����+�������;$Fגb@�	 ��
���s���"o�7/S��ͨ�.>~A�-J �2��?���2ZQk��,����=�a���<�ߥ�N����-c�{��`=m�i�	�[���w/�� �OE�	 \MG/{��r7�/o��f���}���m������wc.ہ�(Y��{�Q�FF?^.��ܶrTp��ebb��P�W�s_⅑y�}�'�Hdd�!j����W� ~#g��ݩG*�?�=�h��˩�r����ş>�}�_�=V)_2�Ҋ\OOc)�p�����oo��ۘ����A���<��5G//;,���!Θh��Ң<�va�����WE��̣$oNjiiAۆ�ڸ�R���{���$k&�=\:r�	7����8<\�ҷ"XEmÜ6@�j�V�0�мx���3R4�I� �z�����f�w�7 �9�Y$�d>_�~
�������RhD7*�#��o�s��Q�)��� ����r{��R����S��:�}镙����mqW�`�l�6;���vA8HF�
뮤�!9.���H`�+]��G3;x�ڳS�Q��(���pn/�[q�e��ޤd>���Jqi*�I]L����L�(q����]lW�������'��A��_LbB|���.ALU� (ћ���j�!�1@'�K��5�BTT�X��������b	�T�*,�i_2}N�nV#�8��N0ɅY���`4���k|n�J>�=����w�\�S��.U[�dK1%9R�jeڡT��|sb�JbӾ/���=Z�����R�f;��eҁ�(�Bd�Ez0��o�,�r��t�Y_8ߊ���wn�
���"Y{��/����
"R�-�Av�6=G���,[7����K�=],������ ���0�5e8.oSy�ק?g4��F)\	�:����6	��;�>�S���W�V���V/���'�HInS ��~�|9JO_���W�)d�?���̓8��X�1A�z��P�8Z_6gQE�N9E3D.3@і���Gٓp�9ts\��$���Y�O���"Ɩa՚l�Fn%%*X~��|�1���{�;�;��n?�,Z�|�W�_��I�j�B�	�v�����+�*-�d*S� F�	��ε�`��w+�m��g���N���c0���em�^ةf�L,����E�.�IT�U&#��f������ў��ש�4b�
��(M�?K��Ą�g�N����͛7�o�q8�J�'f�yN�m�NN_t$Ԅ����M��f����(�<ds��j6���P�2[̔��"D�=oĥe� ��=C����_�����%���A��2����7Eoz}�>HKK����y�MOO#�I~�%�k���[uhM�!u[l0\��_;R��K����&��#Fs��;�!|�߇��v�<:V"�-�"����ڬK9ݭ�E襤���7r_)���d'�_�t��$���*��R<�y�a���������!d��fSㄺ�.DV�+Mm�Ob��<��F��@,�I��xl3{tt��P�4ta��Ȁ[]�++���2C��9v�UL�1#����y�7���K��r�z�����/�K�`m�<]@�@'?���Gf@
�Xm��$���h��(���ț
f�Y���o�ӯ��Yqqq*i��ڥ�Jw�u<��m�DfK%�}���NX�Z>+��y���z���ȃH��+Z����%R	��77'kkk#[[��q`}���$e~]]R��	����"����[�="Ĺp�?;�D�uu� ���뜔Eo����Ï�4�L�s�v������u�ذ [!����9E�C9���@q���\�vz��j
E*�w��GD"eq�W]�gL��o'˒li���"���f?�Ɨ�^~����5׼+V�.�ao�x��"�FP������b�طU�f�s%���(V��i$S4k�����?N���[�^�<׫��˯Xc�l�������oN��q"E�uڷt�|�^3'�@�W�!F/;�I��o��� ��!���.��f����iC-����&��6��:����G�����'�~t��o�E��]e�2wRoD���<Ue�鵘�x��+��V�]�X�g��J�{9��c���$�>G�P	��q.��7�?��u++�,����]��jy�0n�5�VKC�N�l�q�߀;���%�+���c����\g,Ȝ���Ny�y�g��b��(m0��*��2_SBv�?���a=�2�
������+Hi��!��,��-�3��oT�ް�}�iYW��]Wx#������|�H�e��Q%����_��K,�����h������>��9�Z��S��1a�(bbRK���=������L�aO��Fe³���Z���l���ݛ�)n���b=~+�9( �|G��6# �x��w��+e��]����$Χ8v��<�y�������H�TLL2���3����� ���~Kǲj]����������ݞ���>�(��F֣�6���W��Hi#����%�;��rP6��(��1=k�'ȉ�fޝ�Uf;{�@u��^�qM����a���	�I����@k�H����X[�'
؂�|���P�}�9�^�c~��*���Z�`��=��|����ƫ?�}�������u����܆�t�W�Ff������I���&��f9
��-K����0e#�9x���=�{�3�cb�����г��xO=��"�(Cjq�hL�R��+�P��a}6v��S�N*�yg���&uC�	~e)  N���I���#ᶳ�sN�t�e�!�n-��� *7�̈zu�6@�����s�"ʀ�z��P���,`ڀ���z���i�˺�&�xK+�Q͎0�o���'��A�}�@�$�o�0���G�*/dbFzP܀
�5��EE���2�|�z�x�'�%k�Kc�/a-�i{~o�x4�������J�;dpp�pJE��S*�~�r�	�a/����8k�/6l6Ҁ�Af�:E8���ޅ_��_�s�;z2ˍ���5� ��au�B��{@[`&.�y7��"�S����)T��Ǯ���j	'Z&x��L�]0t�A\g��SS�:�.���T:A�	� �%SRO:�<�_⳷�� �{T߈ч7x�#�z��+��������3�&��{u��,������c9�*
L����Au[k��h���G��Ŕ���s��zWW\�t�~�z�ƾ�&l��=Q�+:rr����8���/8�"��ڦՈW[� ೛�7���3J΅|��ώVd��vS����K�t&�u�? ����V~8<uu�u����Xs,W`���9���m`sظ$'�_o�Q"޾�Z<�N�/--ߨ�,g������R��C�x�p�X���f�[q
BD���x�4�ݴ,X�[�ݞ���0;s#�:�X߱A�}��v�^G�U���75����l�����A7Ј?I<&W��
���:����z��(� �c��x�S#Ϧ�Fl�j:�b�<ځ]��u0to�b>�f��!���zns5M|��v�*[���(ɝZ::�?�%׻����xxx�b��C�e�s@)	an�<���\�~��2�~8)���Na!Ҟ\��������h���}��^AE:���R3���4��8_A��萴vr�M�n4(�*��7�ȶkZ�p�$���)�|$r�m$m��%~AFR�Ï\8E�9�]7Y�U���:�џ{��v��
fY������wXXY��`�,U-ՊL���������]��m�\.��#-my���6)1	�Sگ8�l>_bI+ޟjܲ)�����|
�.u3n�ދ����5X=��~��qXFb-b�aʄ	B���mq���6�L��כ���*L�(tc���W�]"w/���?~�$󈧜vƁ�@{�[��6O=��ӻ�|2hSE%E�1�'��"��Ԝ��(��xS�~;����e���Q���x�l{�����Mxv���~D4��\�����_�k��-�S�@�h�i��D��� K�U|������s��Me�s;1���C�i_<yeI��r��>�q���)Jێț^ƻ�~=�N�/��6�}����3q=���[�=�`�!�.��*Ĳē�@'����P=u�s�EV9G��+((���pq�Hz���^�l����)�Y���$o<�]��5f��o�k�;�e�D�;j�S�Km1�m0���[rc��Q���2
�k;�C��^���~Lpg�0�dnn�,��8��H���44Zi��u��U��J����Q{`���Z�p�a�3�]I���`o�n*V�_�"ط�� и�����6Йz�oO �[���=��<�qOy��q�����S_Xh�Y£�H;����H_��j|��_��Ĝ���]YY	�s��A��omP<�!����#0�nQ�v��o���4������!-U�%�������:��}�b�_(7�U�C**h�Â�=���X݌�$����Nd9T%�گ�B"�h��rR�	X�O�ABUC��@'#���� �Kl�`]�v�h����PL�Bm���D����n���OT+�P�C({�����?�A9��upW9�H�2=�䈾G)���{��T�B�� �ł��>Y5n����濟����s��q��|�la�^��A f.���t��t:� ��2���������i�{]q�П(�?�;���ba*����90 �����a����hl���e����3��4�a5`3Ŷ�w�A�QJ��������'a����
`ʱ�+^����W�W=[�����g�

�b聹I��Bgh�C��y6����} ���qɋ'@���WXE������O3�h�F66�a��U�J��5��ܢ����ɒ���QD������L�L�߮;J�:dE�ue�v�5i���;���o�ޖ�b/��߮W�YJ(�=ϯY��tia�>dc�]^���׿w�ji�1�};Y;��VQ�+�^EB��x��D�I_U o��n0���;� {é�OP*R�`�l)Ը�Rc��T���-W:B�pk�ƀ���_@Zk��'�X���vVv��%�WW�Q�[Q��r���`v4ʨ�0ޭ�˔�t�B_�"n{�z��ث�.N�'f�kUc�����
N��֯K��aC���	������4%&&n���)Z�&��N��Ռ��ñ�X�����6��#�\�?���JI1�5�F'��������͍�ܒ����2�.D!�K����E�  �k�f;"�~H���'�kuO�jV�T��ҩ��1�q8?�֘^�ȁq�r����[����a����)�X��+�0�p���<�h �m��{�4�L x�'M^�	[���|��l.|�:�5J�ihb���`-�ӌ9MU��Ý��J ezU) ���|�={���]"��[�|�s7��Z�D��)ݼ�|:܃C;��y�^��^�̋
b�}�X�DY�mE{�sK+���.���=��y��hh�yуҏ�hc��H��ϧ���%���A�u�B��c�.N�m�&͊�	v$��h0דd�DQy�Yy�9��*?��V���?~h::����x�9Xwg۴��Y��Z֣�x,���me%�҉:��E���Warc���Z��9Tr	aOE������w&Ϻ[u���Uc�[�M�rP�r�	�>;�m�2��&�v�7?���$�#��`�_�$�-��V�k4v�X!&�Q�CI�kT����1�%V6���-�(`������ۆFG�Pj�f�	���]�b���âu��>m �{8t�/�3�?'��CŤ p��yг����s_(y�٨R��l��	!]�#�]|}j�����\�{��Xm', G�=�6|��н:��LEђ��EH�`Y<�B���R"Wr�\R���v�K��	@p6 i��3��(�ͽ�>v��0^�3g�,��ѣ �U��ʣ���kk��n�_�F��=~A?V�A�C����uG��p�AS8��;��<Q�f�<�<�P��Z�$~:�<N:-���O{b���zP�K������X���������y����	Rń�
�)�aQ���
�����޽{ ��i�x4��u#�|���g��@R��\���?��o?�^	�&��4�Z�-��ݕ&��q�p�<��Þ�_}��{��7uri�S�>n{����� ���6���D�1V֫�yZ��_� I��Y_� ��ge�Jd��Y�U���X��Į�����Z�X�_���l���?�"9�� �M�w�����O�PN`��'�������T���H��J8iW�P��ԉ�^��4��E������4x{No�	�)~�^�^���� %W7H9l�SbV�J�{?�|�I�Cj/E��{Ɓ"ST����h��D���zR~Iɰ��ڥ��%H��N� ��e|P����%�<��5J�á�&�*mb.q<0�KO��&X��׸�+�$y{{���ߓ�$I.�c��|����@]9���P�Z�Jc��%��K�}�c����>uD_9c���
�J�S~ު1���4�<8�E�v�嵦β ��S�2d�j�� e�d�d�yG�
ٱ�bX���W�g.�F'/j���g>�ty��-�E�~
�o7#����
 �AT�(�@x\��	�S~zz�{�_fS�pCE��Tzf�=h;$��OfųM1f_uѷ�v�7E����� @���xE:��Vx`ǚ����� u23/il�ߙ�
��X��#���Z~�4�4tt��i �GFX��4~2<����Y���Z���߅�^W;�6�.���v~�Gκ�-\SasM��Q�8W(�ĝq�KxC·'�Z��,��~-�gs��,.�\ۻ{hk��q�O�)H��%x�[9�(P�Lm��e����mݑ�T��j��ʄ<Kr��V�u�f*
]޸rV<g����M擛�98�ʣ���YO�٩�u� 1I�#��­TW̣cc�B?��\�*,޶��^nַs<��J�a��3��)d叽�����R՞I��S��㩥�{�2������ԣ�����!H�n����Qe v�OII�n{�`�ܨ`V�iG	�@)ł�M4�͓�������-s���tU����L�0>�ݱ�Εm��x))�����ڙH袠dwyq�k�r�й�[���L�@{u1���mu'I�229�lu���i��D��JY��}��#n�#�N�� 뢾�M;�HG5����E_����~�����Ai,|YJ+B}>�c{����[,|>/bf�O����$=�VP|"�zl��`cﻵu���3��}?�����_�ġ�b2�x���sth�E�\����8~v��$��GB��8T�!�5�e���E6��h����&cɃ��J�M�.�X#o�M��c��5�.V�q~��5��n���|0h��T�n��Lm\Ȝ��2z��F�gt	#����Y��1��8t�����o���k�/�`WV�&W�?>?m^5��� ��z�d���C`>Y3�9��*�W�id���9:�ߋ�����į�����6V�V�+e�M!9�5jt���X����9�?�Ф�����#�ư��7�(	�|��C��xmF�]�ӝ�.�JO71���lMF	2�����T<0nq��U��v�1c�ފ.W߃�����Om��o�Cᡫ֒\��5��VCe� zoYsss�|�+����-��䁻8��4�י�#I�t������z����|�����7���s�e ��Γ'㩱>^�y����C�^E�R���|��C��;�]�i��n�=&e#��HUGǊ�$�x/���㼹�9���e��PW�ω9�9>�ӚG����^����Ο���WĔ�?l����سtgɊ�F_��5�"��L�2��C�ۄ��;�d���Ӄj��Oҿ�bMP\̑�σ�����������v ���Lj�El���4�g� ]d
$d�F������2�K�1L��K�-_��� ����0�3�Nߵ�.�mZ��4�d�\�D>���u����$��xhZ�9�Yİ�+�>����{�NVtT�#I`�������#5���;�ѵ/��ĤY��W9�wV���j�-B1��CQ_��� o�=�s�_C�[�Lt)�Z�4��~����[(5����l� |�Pc:�q���V�apHǸ(�`#'v�9"NF	��u���`�R�N� �:g�E��ho%�����ŷ��z��b��So4�q��IJzM�K��ߦx'W�溱z�����w~��>�����'����d����y�(�~Iy�'��O�]�#5���D�%�{���%A���m~�İ�W{�\����l���A'�tC�0�Io�����0���Ϳ �#6�t
23[T��[Kcn(%����>D���r�p�"��+�2RZ���������!]����7ϟ��@E�q: /���)�?MN^a�q~i�b�R�eveR�kZ��p��8��n5�$O^$�u\V�F�:��d�J
������������뼵[��-���Zͬs�_����|��"G�D}rS����ޱQ�9u��G�����ӠZL���*��|�F��4T뉖��ؖF�����(�
������r�#v�с����LPm7?'�A�ؼ��K��l�>b.��b\���Z�,��� �Ed�v�E@��k�j�LK�fư|��+��E�B,m^��8,��»��j1
JU�;�zj�7�0?��lJ44�)�Y�p��>\V����s�?����u�9T�1�΅*�PlaY4�(T&t$�$��
�^��i�&T���S&RAס^t�^|lo	Uu�^��S�ӊz �!e=7g�R#y����p����7!-EI,��Xq$���Di�'�Y�L���6,7[4cטF w�bXf�å��ӏ�+d�u��;��䰸���'��U�<>����h�):+޵G ����E88�q�� �,��{�Ms�;)�����N��[�C�U9`�{{�Q<�dO�>�^���X�h�OG�VE�H�L�n(�"�,QEq\�z5⩊��~�uu}�V;��1ӹ��A@u���~�����V��}mʠ�zê�ZUk�ݍUjs���]
n�k�75�mU���vě����ĉi���9dco/ #c��AK`�́X�+(���7�q���lv\b�S������܊�A�kV(�@$9�O8m,�5��ݏ�$�����+�+�l/�'J͌���^?]���v�sc��Y�i]� $�)�ݸ	!s�P4�nx)[j�Do��.ه�>\����&P�v�I��K��*�Ҍ�e��e�B0hog��\����L�ih $T��\���y��VJ�q���\�Z,�@��G�x��㣳@��o�F��=06��W�Dr=u�n���6{�bbرf�,ZIac[j�2�������ht��3iQ����� #��W�6��5�u7{8�E����V�7t&�9�mʷ5ǿ�<Q�����]��iLܣ{u��ٳP]T[A!�o4H��� ��Ĳ�ƀ�;������j�t ��3~A[M-�P^f��S �5�>�w�}I�LN�=���P����fck�;�a��q^Hl���>�]���F�`f��|��F8��l���/J���]ۇ�֦�z(���۾�|G4}��BWn��S� ��J51U$f�^��ɇ�����5�|����Y���A
��e$��C�w.Ć\(�&p��L5�ڛ;y��}������,U�/�b93�Qt�8�<H��M.,�� 7����$��S�ZD�NY�O֮���lTgo���D8�$�&�p�ʦ��]?��<�D�#=��UI��`:������F �7��
��<
��x���[UME�Е��2�z���ϟ�⃙ 3��%D�U:
�O��!I��/fgg�k��Jj���������PI��ڏx�i�ڑc=�ު����d��v�B����,$����O����0+�۬,����7��v������{�I�Ц�P�|RX� c��V~���Y�*�3@v�;��2։�"���а�E�XS�	��NBe�Z\���G�E���S���e@�&n8	d�m����������xXa0]_��֖�p��^�K6�%��k��t�"y�N[wߏi���W�{����:j[�L�x�QH���<z#�?E�*�I4��`��q�ߠ�e���}������15��E�g���U�I��nwI�nC�Zӊ#v����{�ɡqzM�OV�;\G�@���*,��QjW���z������(��v)[`��ٵ���t�w �דz���;�M*rkR	ijB�c�Fc}�O�P��0��S��&D(�bf�߼gn��g��W7n��m!����j����D~c����%Q���@�R�|y�t��=ty��{�z4��0$� ����y��(㬹ߜ&���OC3�8��ǝ! WP�����T&q���"��_�� �.��ģ���]#�nH1��v���g����!�@�d	�Bz����$!G�ׯ����':��!qxR��:���)U??q�ۤ��Y~VJ^��bN�����ySq=Q��>�Q�e�2ν)����vpȜUWA�"��u����"�j��]8�;1�Yekn��{W��Z8h�i���! S��kvD�^P�+:�t��F�g$���H2 �:�Dݡ�%t��Ǹs�:�����n�m�GAqq/�Իh[Ԙ���P�C�	d?�K��H$J��PH�"�o�79��]�K�:N?hO�`�S�pPS�N?\�h�]}�^�Xz�����F�v�pO�5��+�l��Y�+��Ȟ��6d4߁]�G�hj�%�9D���][g�z�T����ד�,�̝���ͽ5,��,�ږ-c� _n��Elj>V���P����tu��/��s�HE���=��---
]���HZ��75���.0B�FFŀ�A����������}�~��2���|�}�*�q�)\���}�-��[	 ]K3h�{�����p���ܓ�/Y�+EzVTw����ј�h�T��z� f?M��C���o�.�ņu� !c
��c�GF�0�{w��
��L�L�
-��a~����
���3 ��!W��Ư&aU̙���!l�������M#1a�LF$+v��S�LnE7!!r��J|�V8�e93B/nG~:���P?6N+��U��%0�?�ajCF9��^���y���\�����[
7�O�D$��ȭt������@�҅��C����ᢪ	��F4�_	�9&;++YNNN�i���F	 ����e�� �n�8a1_!af�Rq>�S�R�<���Lx�f��0�5�b���e���B��7�2xɭ��Bwe*�_fMϮ#�U���ʟ�&(��e0��9>9kJՠ.�YE�x.''��ߥ׏�C�uE��SP��Y2jt�~�S(6U7�J��������THv�R��S|��4P/^�nN�Ra.���%��Y�������ʟϋ������֟���88����7�{/ 9�h�m����k�m�o��+�r`����re��5�S����c&?�������Z-����%�=����ȼ>�����/��^���zhh�Âo?b���}��I9u�˃�~��;. �?�'����A}%�b�xJ��+��#ԡ9�I��ݴ)go��d����'��<��P�㥦Y� ~�Dv�{A�G#����Vڵ��y��ݷ]}%_~����l�GpzbK����x�1`�.݅�K� ������֏�L�1h�<�Z���#�x�r�;���l7�WN�.Yz{_9��m�%�2��Pű�[6{}�#*/S��2A�r��X��w�^�-������ȉĿ�:Y	�e	����i��^K�~�۷�l��U���$����:oa�f�
m���R��qR�Ƞf �ݥ���0��|�ug'���'�Β]w�^��.���0����Ǎ� � %C�b�<�{�8m��w)�@�`Re�L������Tg�l�E��&��#�Щ/U�&<`�X#̾5لڅ>�z�j�4Yd�2�N�|6���crXhߺˣ`%��d&'t����.A��5$޷mq��"�/t�!sv��]���i�JWI/5{A��-�⫛�� �۴������������5��0	h��20;�cş�%���k����P�+��h��v7]o~ɍl�c�a��	ǀ4?���5����4��� /�b�6�7���lP����nM`��p;X
o�x�7ܕ����f�����K�n;,l�m<(7؝}7�)YuDZ���ɽ4��e���RdZr��(b[G�8�̈��OE�O�����t%�5��#���c�H@PP�����\;�v�T���ں]��}FX�
��������z>��.A�q^(�y��.�&���7#Y+2���}���Y_�c��r�Jtg��_�\��ߠlo�Mv�����Q�G����/���?mFI�Q�8��=�FH8𝛇GR�����B�|�S���q���á����}l�c����Vb��B�^�\������̭x<�`��g��͑�Ӛ7�A��Hp�!BI3~,E�ѻ*������� ��@�m��=}\�����H�- �'S`���� k��S�^X�.1,����;]����MT��=:�*�=���5�E��.7Ut���.r�XS'�ݍWS��i�E��d����u�T��-��0����{��h�݄-��&�tgi�O�T�ƣOa�P�/{�N<�M��A]���-*�A��	LM�����j0B��
x,�Αdu�zQ��*z��γ�׻q��o��
o,�{k~0�ڸ"�~�w�+�jdz�j40��/:��*}�V?�֞���D���Ȥڽ=r�GrK+�m��91v�G10��������I 7�/?��l{y S
���:hqU'����'є,#^���c�̩g�_�����*^�.*�4��7K�NDA����l�$�k�lq��E@�=�H�(_� g����t����c����h <��4 sZO1z@�	a��EEE��W�**+���Q=��80,�������)�R����n�����,k��T���>-�	%[��G2���Y8����r��<7H��b���5�U��)�k���i���OyHmF��+@Dˮyݜ�Y�����uh��R#��Znnlć=�[�04��wV�����t:Di�[���������<K�?�w>�9��9����5>�A��c�̳����G�Np���p&o�c��_��]�p���	h�wT��\�ؿ&>�ŅQ�_�#@=��KwPEf��r���X�!Y�UQF8�%��=���9����ٶ����N6�=���W_��*�?�	%$�YRD��Ai�X�DB�S�A�C���i��]����"~��^?�����Μ9�yΜy�Wgp���s�Z�}G=��NMv��)��K�J��8J\gt����w/)�o@��g�q��cD�7�&����}e�2�`��W�VHF����Y���k_�?/ѫ�c"V��6������Oę�PR�����,'x��t8e�Q׻��G0�ȫ=d�s�bmOً`JO=0��y�V��oB��=,)�E)Hq�z�IҫH.��d�m�,��hfkcm�}�5��~5!+�����9R���WT� ^��φ���P�����&���	55d�R��tX� E<�|M�����
�w��Ԟ�|z�Ĭ���'"����$�}��뎞�#W�yπ?2��k��������'�ɷ����l]�'Ǆ>S��.�;U$��帉"Sv��VG�|��2�vh�w��ߦ�8��L��w��~�Gt���TW��)����u��++G\Ü��	�@�Q�*�U���;�,=���ja+X�Q�(�(��H�ȹ'�b<����1��'�������D���?�-�T�x9�k'��҄���}i�~Af/C��׶��n�6���Ю�F�y�d��㦔Wb���QW-G�Hs�g�i����<:�Dz���Hs�b���M�Ν��;F���
%2WM��Kݦ T\s�4�$��JZ�~O�Ù��k��5T�ʁ�©�DL�`Cd:W�cc�z�4�2m�t�i˄`/ ��tu��q@g�����<�H�U~����l�x����\5 ��M=#�Nv��,�*`ד���/3)��:zId�z/��i��~}�w,������6%�'����w�1���is��$�uz��.�/P<�ƱLw~��(;;�	�:�v����<�0J�*y|k�\5q��҂l���ד�21�`�K33�mJ�Q��i,%��O�k�-�&��Qrp��ay1$�;���u�/
�gy�M?͇DҦMq����{�!]���[r�3�<��$-\r�*�����pnJ[�`D�Щǥ~����x���{��̓�������h����GR��kv-8�@n�2)�4��uϰO���T��Ȉk�|�S ��'2��O��XܾE!Y;^Kn$����I��f������PWq��M�(萬�� ��ëÊL�����]o��׵rx�l�kc���Hx��m/M^~��M"��w��"����h�Mk���g��N�3�^�Kx�*fR�q�YX�Y�gΝ$틝+{v�~6����� �sC��cWAbx �	tQ��V�p'N�W���ٛ��P4��+l?�(6���n�z�6'5 ��^�]��i-�6�g6�უ��j.8^���\*#>��Ǟ��2�Nֺ�g�m#V����\���ù'���=~��^bXR���a��3_/,(�q�E���'dfV(�ߣH����b7���0�rƈTy{H��B�C�Q.ͼ.P��Sذ�����i��<kn��� VOU�5kt}�U�"J��z�`�\C��а6���eۇ��#���Z��y��,`�-�ef��w1��y����7D�r��o�mt6� Lr���<�s}{�?�3��A���]�i'�fӲ-J"ojWW���҂Z��;��� �`���NJ{k����d�?���Q�XIOBJ��ɞ�K�6(���b��n����[�#,���:�--6�5q�2@�f�jD(��tMhyu���M���� �d�}���*o<�
Xcf�E�L�B��,��������}���#��O>�C
�v:|�g۷�E�� J"\꿧Ֆq��ui�kx�J���5?e��p�;���Qr���-�	���k���+���^Ű��g�F�V�ԧ���)��(9���$`���؆J�L��s�ز'�H568iz�5�{)��̺{������8�����á	���)O�QY�9��6ؕ�`�4[y8�ΒDy3�o%�.��.ץo�b]�^V8��3�:���X�x��V��=�_�|T��xg�WflSě�=�xRte�,��c�o^~�Ggr���X�UJ��}i�;�R��� �N��E"���&h�T�%˩�-�8t���d~�/�`P�r�'%�M,���S��-����B�d��=���az�7������K��]Ǝ�8�f�vP�%.�;$��֜��?W���k���u&˩;扟m�b�&��Z�|^���aeeb��M���4���5�k�`v7R�7<�0._�de����2Q��8
��e�ŭ�6�V	] ��n���B�3*ؾ@{��n(8vcT�B}=�ۯ�x�����˂C��v�5nypK��#l����R�\^yGB��mʻ��^�o�#�؜W�}��掆:Лݕ��Z���[����(4�O��F8�Ngtj�8B�bn��2��Z�xM@���� ��3�t�,H%'^{���駗������mm�S���4�ͪ��F_�?wl�j����ޑ5c�0��O�7g�_��u�<�]7Z��;��bз�b������VC�O�����.�������0Ei�5}���t��w7���|�qά*����ő���+�<�~A<e=l5Z��^����K���^��g�r��b�9�M��g�
����}pbPߟ�?%j�Os<�
�(��L�di��E���3��؏�Bஓ��l�T�,F}2a���!�_���/�ȫ�R]ΒC���N6%a��G�����I
���w�XHC��� *;"�:;�i>����+6�ʻq�:`�9]Դ�=4އM���j������'sU-!]ָ�f���K��5���Qؽ���@������!0�C5f�m��ڦ�Z�C��SS��o�ѝ�(�����+�Hkf����	��)���x��^�6���nd&}/�������I��I���pv��V`r?�aJT�0�����W{;�-�;�c��
���q��'��<�rO�e�rUMH�'kr�T���^�%����Ǐ��Q��A�.�?�Q���Յ���gs��ܕ6
��H�KP�c�:n͜X�͉����x�����Z�f���Lja����9�����o����sF����=خ��Jy�e׹<?,������ő�A�1F��џ�����~[ݦ0��C�D ��6Lc��#��X����j1r� !1�Wo@邏����ݚ�y]��/Vŕ[9v���dӥͨK�ww	�����U~�I1�P����j��7�Q�x�S:�̐�7�r!����'ۤ����n�ov��	��*&7�T�d��2#����{�Ħ���nX2��0CI�R}0ť�k�O+�Z��,L����V�%�;�R��-���SL3эv&���R�V��J���(��:�w<��E킻m,�y��-���Z��C�7'��s��p㏵���>Ϣ�9X��d	�0�)��&�
M񮷱�ǒ�I@ۑX�KXԌ`BeJ�����.^�Ձ.rO���L��,�}%k3vύ��+��Ϧ7�w��OT��P4�I�.5������>4�2��Sڤ��[l�:<K����uK�kc�Y;n�u{R\���md݅Gs1sb�d,�6l	��:��U�{��
5�תTT!�'���,�m���B����5��-�C!u�/��=���4�����mK�_�<.�*M���f��.`�iƱ��K-#*����y��3LN����~���9&n�X�9J������O5���E��4>��By6\��N �r���SѢLq_��]cl`w��Vz##{�����	'�=�a��;���]{���#V�TA�,�W���1���L^	E�K'���0��`:��.�:P�ۧ�P�~,s���\�b�~�w:o����-���q��w0�^H���s�^~��:jb�^�?
�h���V��0c�lBccF���g����柜S�w���&l��z�(��g]���8�T��i=5�O���V��zs�?�t6/��Ll��<�'3����A8�<j�k<�d�ږV��u�l�.�4tV�(Z'̎I�_��>�8������,��K��vv.8!nu-970��eom��e� \L�$nP*r��(�`9i��i�q|y���N�����Z��u���'/	r �;jT4�R���i�K��G Ŧ��o�R,�Y���
�G��"�nb����N��o�̓�i�,+����>�Y2�Y�6	�)�u'X��@	w�� trp(^
aX��c������u�Z~�L��ҭ�t@������;�n�yiDl��l��6
���}� Bu��(ؾfS�c2�~E@������:�#��kyq�`qK-l�_P���������3��<r���Y::�~�o�p�kQ?
�<�S��<����W��wF���|�B�7[�:���1���!��#[�0|-�\�kv$EL˥99�&
���CT�j4�)B��+���7��^u���#C�3���6Y���R�e.ڟ�l���d��>�ĺ� 
����Y�(`����J��ݞH������:�Ɇ>�D�2w"�VEf��R��ѫWG�'�8&?�B�.=>v:���ȑ�i��ƻ�Z�S����v��m�c4����N��{�<S����N��y*?�9�G86�`ѻ �B ^Ƿ�@5Ns�5~h��V���=	�*|�O�Ǔ�w�(�z|@�Ǜ�rP��[{e�88�B	��s�0
�{���Z8Q�Q��$V7U�N,0.(��}�v'_���d�ϲ-g������kj�-��g��������}�.�V�\����bN.s%�Ae��)�F:���%�m5fkKo�'Hu�{�~1zZOU;vL�A��Y��p�|�P��fs%����Ǽ�|x�נ�Noo���Wh�������S�8�j�|��00�	xy
�'*�g��Iw����	���@�����ox��uQ�1�ۇRL���cP�����zܳē�5ν*@���� �.v+'2�/����.�)*�vh����Ǿ�j��d������_�ƫ	$��p�e�V���.�a��rP>�T4�ш*����!"���|��F}ҝ�Zş�������^��RXq}��R�zE"<�Ok�/��f=��⮗�������#��X�M㧺zn̜�h�U��c3kȠ�*R��x��Pt�$N�����/ⶌ��]�ё�[�I69T�nc_�p͉y��	Ji�ȋ��_�0�>W4�ւ�u.@G�`��4�3�E�r�3Q�T-v��'�%�g`��ݮaN���6����+�#�c]Z�Z!9�&��@X�bHhi��$K��}{E��U�B����6)���.��>����n^�s����k�����R�D�c�7��&j���D
N�����^VC�:�
�F��O��^�8�X��]%�0�I��n����w�ݓ�p�Q����
*�b�4�[���Ӝ��YSD�'��+Z��kQ��*��R�y�" �����
"Ï�{&�W��湄��V�.�@����	R"TK�zb���QP����7�� �^��j�G���Z�LG��Qou~����߉h�">�I���C��/�w��*������� $tO�]�P��^��<%��� egHć�É���}c��<�(:��#�R�}D(���HA���ø�_�~���3P귦�XR��g�{��Y����������-�*C�w��"	K���T�ˉ�� �>!��N\���f��3��s~.�-~�(a}�"��ܚ��^B���<��		���)��r�����~��Þ�~ s�� 8j�	Q���;v�6��"���y�zOzWl�-���&��]��>��1D�[$6�܌JR�<`+s��<[)�W�G�\C4����;ܫxe*{��fl���%H��;|���A4~&���,li�qC��ظ�n���tje2vf樾8�a������ɡ?F��|W�kȓ���h��6�ũ;&�	�H���~���Vj��k}=z�y��/ʷ�2}�J�'t��	Ҟ{ T�0����>0��M��|�G�~�~�mP�-k���g+C��BƫR�ǧmyy]�o�{��m�Qeh�z��Oa���V��jxP����r�Z;������ܕ���OEo�uqWS@�3�A{�H����8sFs)Om$�/��aT�;/o�������c�#����JL��c����P	��ZsqeI����Ζ�Aa����b�w���(��=�D1!أd
ʇ&�-��/r�k+�[<��G��TM�n��zG�Z#p��+A�6n-ѫ%������Ye����<C��T)���w��E{�� ɓ��� �Iu���É�XV����J��l�٬���Kq���/��E���]	t�('c��7�kbYY5@Լ|劢�`���܎���î����Ù��iaiJiB��Qv><���wG�Lc@�0s�t�%Aۃ� ���/���Er]"u˘��]��}�S��U��V:y��g�w
-'�ߗ�R`l�om�ޡ��8���F���Rt����)L}�+HLCU5
��ad4��J
���?d3tLș���#�f(���k�N���أ���>W�12\١���3��O�g���qU��<�]7t�\�H_�J���U���z���t����G߇=x w#��H�6O���+L���m=<���o߳rU�>R^~����nM�u3n)h4ZA��5�9�*���&�m��]�腕'���h�Ј��C^aᒑ5������li��;	�6�;�9Ɖd`����)�s5oY��q׮�}PN�M�z*�!�E�Of9����N�:
+�����L�-����=� 8Ȅjk.K- ����r�󊒲������h�-G���6KY��O�~�U~iV�C�?�B�Gg�[K��W����S��,J|��ɑ��i��\�o�B��{'=nyyy�LSUُNp��3!L��/fc���a��n�Xm��ɋ0V)�8.�XX�s�)�^W�tI�q��ɸ]}43K���G��aBhhF�n������b��R�wC���c?��񂢢e�-"�]X���|�Qt3��8��F�n��{�<s���f�s>�l'H��>f���ي���Qܽ�M�vV�rg<�I$�֝HZ��p������b��a,qrޤ�x{�o\7��ɍ�8�ʠ�zX��V����@���g��_ۻkB+LC�}��|��� s�Y�5[����lvCL��R�wY�����o��������$v %I��ξ��.G?:\h=rFID#Z��	����5���h�"ǎ�f�:(|��w�����Lpf���-}ym����\��`I	ｵGT�z���[ʗEm����pd��[��[�X�c���ǿ�w��������5��&�^�NY�SR�n\:���>%W����^t�w�(+5}��13#�(tFݪe�;��u��p���sؔH��KqCXņլPW�"��.EÏ�����?�%Ɩ}�l�����*�R�Oxdf��'��"��>K,���|<�.�|Lom=�
�
q�>���{(��7>���Ւ�m�(@9�v�Ѷ�.\�O2�u�/}���p*��垞�V�N���Y����/�O��ygy�z\3^�f\�_�G�O4e\�t�n�3�j8h��C#M���;�̥D�NR�A�6���YJ<^���|�	gTE|vS,�E��.��$���m3���~e��W��/m%���c~�VlCH'�� ���6�t����Bŗ�$aVy�阯9|�%P8�������B��1Y^����rD�T��FN�
�����.�ܷ���1�mz��I'>&��<�5�t�\��`�ݗܬWՓm+�f��+Ԛ!4�7�W��s�챠5��o� 4��]�`���-~�n\�ck��dm��Jt�j0��HEl��a���0gݶA��_Wf�0������u�������X��b�2:^�~~��h#�^�x1D��L�&�����C�PX���b3j���A�ռ��Pw�aig�z!L�06�Z��r�5i���)2sJT�����ntF�����C��ABy��bܖI�<_���<�zM߳C�c��E8b��i�:$�!y�Dv��[���+�6ϖ��t��ᦄ���Y��'XE�aS��o�M���f��� Cfk�w�K���jb���WQ����X���܉pqM�_���y�@Xm��
���H��{�$��x�N`lF,S�z�=���/lmG�S�>_H�TU�_>n��z���I~Dp%�.a6GKm��5��m��HɆ_���K�o��P��>11"r�e�s%"9I��t�i������&�ΰ%�a&-͖�%k�m�ǎ������Y��/ x=��႘�='a���Ld���\���EȺ7"P����"���?�=��=��-:�Kg�^��6���9^���m2F�o��P8��\�+';XtI�Û��^��:�Yg��%���M�j�m�g���8�I	6���9X���s�2N��o�B�Q�����ņ���m*���覾�HHI��et��ɍHs��>�suB����vRc3�n�;f_�#��͔\«�jkD�ˊ�������V<E�06�.�$B:)��F}~�3�4E����P�b�;#cc�K8�h�tS�@Y�(����-�,7���jg�t����N"�9I�׷�7���z��b�S5\�ss�a��ϼim�q��bB�K��\n���.�fU��O�U��s4q�bk�,}�� .֞P���L�˯[�:�e�8�m���Vz�ڣ=�F���qA�?h���7~���iC��W��O�B5����R�*���S����`��NNN��ЛU���x�f��l�� ߤ%�	zH��z�ߧy��p���M�j!֢?1sm�L��'*q�{EO��f)n��x��S9?��C�S��3�z��Fw0oZz��.�(�W��i	x��s��=k��i��basG��q "M9��Tۄ�%'S��U,�ޅmz@����k���cd+++!������r��pg��U�T8�_��B"�p�'�q�O���iٛ���`kr���$�I�0�	>{5���yG����nN\��/�3O�k��}@��D[��\=��V��S�G)Vr�Y�����C��'�[� �O�J�Btnmo�<�]�V��N$jiO�>�w�S1�3�q�Z��Ҵ��quY�:�K�zl�����{sAK��˼#7��9s23O�9h�F��ϵ��ׂѢ�P���7ta�7q�o3�N�3������{��ш�΋����FX੣k��)����M�ou��E�S/�F)��A"K�
-Ặ|)��IC�`|j��,���Bֵ�A�W��d�b-�W� AĖ_�M��>s.��RF�`9�Z��,L���ԯ�h��z�r�=Tkn7�:�fz+�6X��������4�'z��8�A�y����R�������ZҟN''�� �*<$��#rn��*����Z���(�<�H�l�iC�9�J����Ӹ���u������3�13�4>=�y�q��5)�^��Ɋ?X�!��0HV�>����/��gff�R|��K�M&�ʃ��\]G�L)ޣ�i�=,	�=�2=��J���0!��p\�W^؞�V��Gv"0[8q��`^@��L-�#���.�@�_��'�����\e�2]H�a�O����h���4���]��څdK�:�T^��ƍ�vḷCB�/2�E�-��i���y�ڛ;-*��p1{����455��J���>j���`��~�*$����Q��P����K8cw�JY#[0B�K���o�fjj��y�<��P-^�1���f��$'��^&ك�!��V�G���8�GGW����o���� %��-9��oO�a�"�8��|��+��~�
?��@2ZV����b����]��Ǜ�K+]_�XX�>����L�އ��^�*]��Hf�����GvrQ2���T1�$dd}�u~����/�s�=��Z@Vp�%.#��l��T��=8����FIB�p�{��f*T;�Y�r{�F���ж֔c7i�2��[�̈́R.&�i)Vƚ^�~~0.�\P��|��?o����"�ǧOuс�z�2	|[>tpS����:���0/O��y+$k8�*�˷o���-�$t�s{���A�7�B�[�=ys ���r;��p�����]t�l���D���AK�ї�M�hƪ�܀6JEZ:(9%z[�?����n�Zؚb���D>��塳y �ڮŦ8!��p���\���I+P��h[���>�8�`3�q�W�aդ$��͖�	}ʜ����=����o�)4����_��g����\ޝv�^ꍃ����F�i��+���I�^��C}��
�l�xxV�+^���|Ms$Nf��;t�0�Y��=ٞZ���;/8/�q�4��s��B��Ѕ�<��&��G���џmMCC�񵍍��b��,���Sر"������nk�3}�t�.zh��4(N;������]\�=�$���ƥ��M���6ڊ��\�j��{Ez��nk��KC�������<���x:�q�}G 0:�v�Q�$�j�B���� )��=7D���Y���rr̦˚,��h�:<^pP؄��v`6V�#�y)�r}�w�h�M��M�I $EI~���X�,��<t UP"װ4f1VRu��pJA�u�wy�V2�a�����}x�@�
�C�x�Q4�#�lS>�_�y�M���Y^�m2ҧg��$���=e���Ҁ�i������>�H$�-1�G�g�x�"��d2�\yۓX7�FgA�S�hFS[;?�۲��^��Tyv������������������Ʉmmlz����f_����[���+��a'k��w�@�E��=}�i��s5P��6L�8:2µL���B�cR]+`Rj��5�����D|�m��|ĹYF,%�`/�n���.N����j����#~�Ït����j����Q��P���2  @�.�����5����bv
	郍�;4�������¦t"}���|�0xX�8;'���Tk�>*�?�9^�˚���Wv!�,^���r�O^\)�·�pB����R���xyye�5TT>|������`x�T,�A[|��"~���+�:88 �&R��HPP��q��w+ ��PȯN�\�r�x�W�{������˭**-龫/8�wl��0�T���Nc������{��> �斖�YY�G(Mwwʘù�֬�����+<|��m^��	0?5� z 4(((F��0��2� ZW(!��AZݲI/_��  С�p����T�|�j4ONm-X��Җg�>�	~���Rmk�4�*k��b�W:E3<��1�l������<����o�Ù����˵��F:��@���������u0�ɤG�oO��N�'&&�E6�#D�R�������|"[��'�hьA�S�R�t�V�*�	.���謯ܤ^4���N[���؞iG���a�~(ƅ��s�n�����)Վ�낪��u��	������W���V���!�[>��L�������ܐ|��+!��ɩ)H�D��l�ܬ,�P2�1�wJ�_'��`1�j�	�x]n���N��&9�q���f.bv+�+���J{���5μ���S*��0�ȅ3��ӻƣ[5{o�9"9'8���WwY���B�%H�LSCC���<��3�+4>��Lօ �������1wr�A�:�Y��pk���?E��M��f�=����1HU�d9y�����n�S�߿�=�&f�U 8~YP�Ch#����H
}F�}�x�2֔��	D�6���|"�{)��o�����o�
���<���F0�еsx�5�3�w�xl���n!t��1�萸��CoŇ���څ���K|^5�
l��AQvvZ�N������'<gJ-iY=��;� ��yKO#���[�Y8���RfK����'þ���%]�w�mf��o�y����쑑�3'8�H��^���g7|�͙���4��(5�Q#�^���yy�G�:��d:��{�	�*E0�6��{�K0v�#sw�_�w��;/�d�z��`"��Ar�V�h$3m~�
SN��a�xG�-��uHIz�'s݂��2zO��^Hɇe6� ��3�c�{H8{~�Y�B��|D! �*gP�<F�5��{_j���8�@����"P2A6�bֹ�,��5�b�|iVś��[pB��Qr�'�27���7*��uT4{O
�D�x���ɕ��6�'�c��� ���g��qr��C+�(OH��mʎY���&4���%M>����d��j�WiE���K
�.S�7��PL���8��ۇ��[�gZ��n��1�����·wh��:��������L�P��o�3��� �ܫ����;�b�;�Mי���n����O3�������&��N�y�)���}��^l:Q�W��$Z+/D� ���ޤ 9�ΪO���}xi��ۺߢ�������h�x�}�RF�/��9>�[��?�4��C=�S�p���4�-��܆pX���n��/���DŦ�:Ăg���� zB�����TXJBHq�_@V�*Z��[Zyj�3E��vDw�Ŧ��G �z�r{j`�g��-��%�-���\W�w&���Ҁ�8���Cwg�#B�3�Y~�)�r��|f?�����O˴)�������{� ��P�T�Ҕ�m�ȡbO�X�z/R�b��c��{ͤ?�Z�h4����>���}}U`4�6W��j`�TU��;9>,=��� G/n��T���`�`�]Q�Ң�3�Z��4s����������������!����|�~�Ը�˂���{ISM-z�e����q{PH��ȌR�`����g����PN0�L(�~jo_1-��u�ζ��;~GC��#!Ε;7iJG2J��ˑN&�Saa�3�]�c�w������82��BK����Oթ����9���h��p���.�l[7�>���x�ծ��55Hq���+ �iH�5 yBK^�up���g���FZZ�P�"Y��E�'l5�j%a��c�����fݿ��Pڎ��"}'1$֢ݺE������72�����n�ś9�>�>�i8��B���
�e�"@	�hޮ�c�vT�k*���u��,߇�f��L�$�1�s�!�����=j�[�L^�7V�Q�J ����É|�Sk���g�����6:��(ࣷ�{�����g|�����\ /���K;��AK�zz�9#,�& ��.g��Чb^�$,թ�%e��I'�.��ׯq�0� )���s�K	dx]�U��폊)�D���R�;��h��^^��~��HG�F������V�X$ �ɏBUD7�A	F��R�	>@�x6}�����z���m�N\
|�ZWp"ɡ���I��E3)rH���W��g|����!� 9?�6������cc�%i��Hȳ���X��>�ՅG��]�����\Qy�z$W�Sr���#b�Y��V�L}��B����U�=$N�/K#�(I�n�mC����>$���k����Sy����ݫ
����--/�]2Ժ;� uK�������@|��zRq9MM5LJ�v�I�{oM��C�ZQY��VId��rv3�� �U�.G����qn����,n���C1���抉$���W�N�:hoA*��47OC7ůj֭�5�E�����'_�ЕRv��)�#X���-W��p�꺦l��[
��/%�`�ia#ԣQ{����Wu�e��J�p��MRR��!��'��V7m��CR3�G\����@X���[�>���O���SW`U��t�<�xX���tX�+,���MHD96�GŰ�[�� Ń'�L�����J�nd�D�ýX�H/\�
�~+�~[]�s�[���j�B~F�OD�逸��؊�ȓ?�lY�ᲃq成�=Qmy�/s�����55N:)w�B��yvW͌��z�vc�4Q�H��#iI'��5A�Z�W�6��{��L�.��U@�+'�ٛ���k�Fw��+�T�(@	b���9#T��f�/M�j{��*Z���������,=��ګI��P=���H�*���Z���f˓��^��_t�F��с�d��?�k~�h�<)ɋ�ia9,y�%S֮������n�m���u>��zӆ��R8Ru���1��3�)&d�~���Ց�[y���6�����{.3�je�V�}�|��@ ���k�B�5�r_��ӧ�HU���谸�S�7ɒ*����A��|M���k_:%"%�A~��6���ǈ��V��~[��N�&��Z��KIY.ˋ�k�'��Y�o���wp�@��ېB��x�8[_��q� �S���2���.�4����2w�p�f1��E�?KȪ��\ֲ�WS]��J��)WO�^oH��W����o'��V×��h�x ��lû�-{�{��}^��5�$�6�V����-|��q�(C�#gs"e����o�ΕΫ���s>���Eތ����%��d�G8<sg1����ߺs��b��e;C�����g�m~�j��ϬpR���4��<Djb�l�)6.n�~') ���]�-�G�����9�#XU�ü� �� %�����*��Z�\P�
���%�r�K����z@�v.h�`YYb�5�W�:sM���8[uL���"�#��B�V��}�!"�����?��������N���NM��a�Z�c�bM��]/��STbr�g-�2Q�:�{_m[��s+�s���+�4n"-uDq~�4�E�7��Tv�[[�ɼ�|)����1S�u�V�B�74��N�h���v���Y|`���q�u��[��"��᪓)��	S��0�{?��m��r��T#Z:�]��z�V%�����%^��}:�^��l�g�[ib\�D�֞Z���3���U!��.	6m�����Yݔ����ann^x��r�*����$��%���J�C�q,�E��FJ���BVn�S!�u��M(�FN8��o��[��9��؞H�#��O�w��Kr��٠�(���������R���((\	� ;5�R��3f!�JW^�ܸ�-�wj��-�g0+Gj�٪��ܠ<��`L�=�����A�D�%R3Ud��贺��)����@�3&�;��_��]>[�\?q�r�~�~�":Q��&J��A����t��=�q���jW){�zM�]���#:{��ʩ�!C�"��",�L%�w{{�f�k����l;@��F�����S9zH�h�uCBBx\�@\赨�����E[��\�9�[4�<x� ��{C�t!C����}��P;M�'֭�  3x���?;CtPf�ȟǓ^�(��7�w��W�|���w��t%�c��Q0��U��Ǵn���+�@�ͭ�/��;��}h�c&��v>��s!���4��M�s��	G)�e���iJ���ŵ�Z���1[C��F�K$g���.�1k�wx4��:h�`�=�m��ϳ���������U*c5��E8�4�w0�~�Q�L�a¸����� ?�b�t��a��j )��H��y3����
�-OʭƵ�,�EY�rɗ�
w�Z��5J�O�I�]�W4(m��ߺ=k��d8Fj�f����-*(Pn_�D'3=� K���4�I���u�\�����ESO���:@J�g�A�����:r�r��S��j�\�� 1�#�]Si�}���rߏӿe��K�y�t~����omu��^o���/��j��pPm�H��g����J�82�ͫ(̜�۫	[��)?5�l����%�Yk%g��j����ݴ|��{p";�O����f��8[gТ�0'G�]mE����qtf�t}�8����J��xxx��Uuu� �_��������ԧj��zL�|/2���}���>�&x5��sZ�W�B�g�}����O�EY=t�J6#���s�n���V�|�CF!�����Hq���.@*n�c�*��	ZliY7Y{�_H��|�x�ޔ�ib�eV��bI��N��M93#�4� �� _�1����mw�ɇ��._��#,|����m5!P�㘸�u�񜝝c�A�\Z\챐���K�11�tn�_�@��Q�!Y?o�����N�z����bS��6�[�ko��+��+���k�����Ma|�������R��O=�"��v��b��t�;�.,򮟚}�/1O��i�~zg$(���
Y�pG;XR�=����zT�}��Znn{SJ�=��q=PM9��!��'���	S�x�5c_�p�B|ݺ��
*���v=&������H�"yϨ��Fad!buX�{wb[��������@����?_0l��*����/Ūԉ9�?�ȋ�����H����o���Y*�*ٹ#���d��K��W�eo%t�{��$f�\���>��&+'l�<����ˬ�f`���q��/zc��G�cr��( �ⳟ.��Yg�-�&�ȩ��x5+Ñ����_i��)0���̾T'��%��'�[F���\�|��R�j�M���9��kcE����:����8�W/�����#�F��f�llj*=�Go.go��u#�q��qO=Pj��˻m~��r99��&�&�9=M���% "��vkE+N;o�|�=�ƴ��ѷ~s�uI���8�Ie��v. ���D�d��)�d��P������$�l��R���T��|�=��:���Z�^X�%���������{ID� W�����D���z����:����;Ϥ�v��zՊ�
�������n�Ր���������_pI��i����w(R0p+=]g����xJ��ԟ9�(�;g����Od#���{��d��W�H��t�=���"> �tʲ�_G=��r[myQ�]��[�����I��b>��N?q)~?������W�!��&���i}���7��p�w
cd�ǔ.U9���*X�B1�,�r�(�/{{PH�M���$m��*>d	�Pa�i���EU*�դԫI�S��:LW�,1����pÊY�0ӂ�o�o�D�6��>�S�@�GSsq�r��O� �͍'��H��W�͠^e��}&1�fP��ROdr�.�?��3�Ҁ:��Qq^�z��\q�S��r3o���25�c�wT�M$s����-�I�����M��v1��l��]�fKL.�֬K�e��O�A�d�����8�w` :������p�y4�������[��]�e�oO6�Y�҃fo�|�+��~�����/�2�r�(5TF[_|P��h��oб���� ��Qx�H1߃��N�>kk�DD�z/{7��Z[�K�+�m����� ��ׇ�6��"��p��
}ZyY��
)[�B�`�;���9�~���d���2��D8_�<Q=�bX��O�0��X�9��o?q} � z��!&�L��O�	U.@	�g��z�p	��,˙D���|7�n�'@��oD��x�x�ߝ�ŉ�ɯ�g�m��|�q�����g�����{;���U����8�jF	�"���1��U
�V���:Y'�pg�'�D�~U���=m~��}]�SȧUp��n�V�����¬��������۷H���]$�e�ꫝq���"L�=J��Jt�D��oD� �UL�{���h ܇�6��R�MW�5���o��y�*I;Y�Ք������N;���������mJp9>����`����<�
��3�v!�0n�n�1/��'��n�?̽wTT˶=�r�k��((�@R$K��Ar��AA���dԣ�( 9#H�"9�"Z�d����n~U��w����c����Uk�5�\k�]���x�A��F0?���B?��p�>%!���l�TE׈�l�^��w��*�!v��/�6��@q�x��}]xw-��Z��wD�X��^�#�$��CO]ͮx�H|⹚�_�_�N��G\�9K=�2�Cɦ�;s/�6��ͅ/�T��:�,ѷ�@K8&:w��yI�K�G��Sƣe	LS33e�F@(e����Xo�D��aUS�/����y�Ƈ��>ݍ�vA��?ٳ83??�� �Bl��+m�'��(v>�cYI'�>넫��:���������o` n���m�[/�T��v�\��:����Ļ}�W��d?��J!+����,Z�ru���͒��tW��N0D<̱,���M����������u2?�jxs��*������/��l3��O�b�e��(P��� J�jLM`��S%f�����:�P�^����ss+��iQ�� )�]���}2>z��9
6#y6�d����+��rkuOx���.6�\,ML����%#|�������
�����率cF�l�f���5��?��?�@���L�@.�X�@�y�ϕ�E��X�R����N�����Em��H�2ӹ�Wh�����E�N�P�����q������.{Q��1����̹'@��DK�����+��P�%���;]9���m��h����8�m��ҋ���n�i)-u�Y ��#t�G�<��e�)_֋�ݹψ��_����U���o��>��i^�ւ�m\��[���y�"�r�bq9�gMS���6�e_���kfq�,�ZMEW7��������)P6�e�����,�)SC��%�Ǔ�M��V*��P�;e7�[���!wsn:������ Ǘs�"g�/F�pk�GN����Ѱ��܎�:w���k����K'�*����pD��<��s2a�;�\�4�ǌ^�{W%'�΢]ԸjC��e5����6�4M���:4����^߄������O�|ic�RK��
�ԩ��\v^6���JkJ9�|yp%�X�3!;�p����M"���2P��I�	���j���7a��}EEG�����{�d}�#-2��0F�P-��סɮ����o�Ē�i���ܻ f8* ����l�TW�v�-g=����d�h7�Ժd�uG�����)Ij�/�1�^�>���j0,9o�ol�b�������%$��� {���T߀�.�=� G���A8�Q�%>�C��z�0����vVU����s�t��IU?�^��cf@a�I�bw�Yh<�l���,���#mˢ?v��7M&��w�R�.ix��J
nR��(������Y��*v!bJ����� �Žk�Ϋ(����ɮ���3Wڽ?�)��P��В�t��/\5���m� �M_��8E��u�1�
HZ�'{k�r��1Z6���:	Ӓ���9���H��$�p ����`��ͅ~�P�kxO�2�7p[�y�9m���FZMx�w? ��� ��fX�$M����则�%n=$�ifu��<@���Y�It������S'��' �̞,��u���"~���Q����M��@�uC��d��%Jȭ(F���@K��/ϰ��" �R��h2Y����=bt��i|>Q�?Rb_)\��q�HX�e}��V�9��=�<|W8jK�WJFO��=���wY���󻒽ڈՊԸۼ�_�� .��G��%�:
��BPb�1��=O�Qb>I��^_�$a�����B�*�%��5�P���� ;�\��-��m��l���L�g�m�yl�������|�`���j��w�J^NAa
����]Y�?.����\Jg�v_,�4R�Tz���eY4��p_��$�E+�~0ӕS͠9����лsYEL�91�`|n`��6h���a��w�a�+��Z�!c�a�5���ko-�.+�8�C%P9�Y-l��[]F��O�I^{���oE��=���=��#.����M�
6`�>~�����#J�N�_R�yY7n���;��2~���'K3��qN��*u������)G�4�^���_7��z���I��iX2�L��败�6󰓛z���P|�?��=��Ih�s�k�-�3I$�rt��ٹ3�!fbWt��+�@QX������W�
klL������4�����k$�.���T@����5�%�󿠷%��:��9y��O������Y��T������YRT�w�Ц&� A�������nf��Ѵ9*W���>|a`+ۙ���^�p�w������3�?�� �dV'�|Da�В�yN�4ũ��^���7�	�#h�33i�߾�
����o���_�˺/!��ٙ8�0?�,Mw���MN��{���7�B��f��p|���s�(��C���v�$]S��폯���J���+�h�}=�%c=7 �j�;r%�A�N-!+���p���uⱚuC�]s�!i�T���d��ﴪ�HR�×o?iK=Q:�DԖ&/o�D@����l��\�2]�X �'7(�ϱw�_?DOFi�&(>U�ϟ%�5ʗ�l��ګ�,@X<�Պ����j#�hy�w�O>�}8��C��V%���<�p!&fT��fc��-)��d|�� '"������tUDk�7k��G����E!�MP��N2HX]]]xC����P�~}:44�Ɋ��_9�2|�f��M���B.4��l�_�$,�72����Б����Z�Ί����8>{Y�u�
�������8K+����7\� � ,,V�;�y:���^gC���$����a�׾m����O /������Ve���_o��7���}����.���ٳ&������j��/nݺoUT�[DF�^�SQ]=�_@ �+E�[5��0 ��ֲ�3�]-B�Y�fX��@(l2��×�̯$�����_�̨07*��y�g���G�V�\����C����k�'){�>3�-@%-�f��W���7v���$���{��{�y#�51��a����� qS����|ޏ<��D�b@���%�g@Ut篻Tj��� ��KYk����Q55M?}�̤���4n��5���˵�/#h4�$�d3���v#���9e����̛�Y�~��v����j�+�� �͇��y,\�����Z��q�Vgg�6J�(֍�~���J��OJ��=�]��O���]�_�y�V�߶IXX�9Nvw��,�u5��?�d����)G ��[�����YwJ*��89���a������gώONL01���O���^�Z=���鱍����j}�ؾL^|��ӗ�i>�T�V�	&]	��_���%�̌8-#��P�0�{��&yy�����.{�ؗ���%W��b����v��Qa���gy�$tt��'jS����N�f:����.���?(������/����3δ� �g�u'p���� ��D|�y��_�����
h����R�W:l������E^3̋���#�s/�[�>��#���0�;��AeZc��R�֞��ӎ;��yP#lV����%UgX��Ek�t�H��y��iǙ!>C~��n���B�6${m�LF�,��R���]��j2w��,*3�6�S�GmZ�LI�yN�+���#�a��Q�@�r�x8��L�@���E����ٷ���a�pྖI%�p۔+�]`�cY�?7��ͯ��;�ę7"�iߘ"W��xO,�|t}�X�!��=��ä�@��k{D�mS�=�ϯVj��?���􃅦�i=K%�=�y_��	m���xVN��S�D=��k��oz`�Z{|T�l@@�٨�{��֩õ��Y�.UѝS����S*.�Ʊ
-������H;����O�j��_��U�.nx
3h�0�$�ŗ:�?��sw#������v�����5��6��EI7�� �1>K�����N��=>N�mf�JBs����6P���CC>����g�Z�s:���5��{�d����ș�S7����k�Hw�E��)L�������������
��㧆KSt���\���F���{��9=�"���}P� �V��~ġ��:�I+5�a�t���p�~�
Bܾ�)��5��a�Jfq�H�y����6.�&tͶ��Z�!L��~cᑪ��yw�d��A�o�(����z@��rI�CkI�J��& %'0nX�=	�;dx�*��wdj�/礇�VrS2j�?I�F�[�T�Q5�Q��}w�>�1��U�͹G�0�����JUQ�y��ǮX.��9;[֒��:�?�X᜿bk�E7���f��.�y�Z-��b�{/�<��S9]~�2����U����?{YԻg_�p�X]�֘���z�?�m�ֺ_`�^��s��SY 6�±��]�]v���qR��o< y�H�".����C`7�2xL=�0}G�Y����lN!�x��믤e�$�����!�^����������~7%����"�9���fJ�'e�bw����9]�ޣ�O,��]��Umc;����$u��L՟�+���ā�68޴��`�H��)>!ԡK�v�◦@0JSu{Q	�{���J�;�}�;�P�����ÙQᵊ�z�iXt��՝�ϝ��)o���0�>�!񘆆�������Z�z�h�<G/�uu�Bf�cL��>�,i�\K�ұ���'��6��ǖ�-�4�?���lZ�"^�\"��W�1p�A�y��T�,������W&`� �\Y�l��$	FjA Wa�U�p�3��L�|�}я��^�R�?+ş��i��7l��B�������d��4��mw<��{ש��s�ب����J�(�����f������v<�R֖�p����F�bt�v[�ZӴ�uWBG�f���@'.�n��y���N�|���?`���wс��ן����D[a�co�֑��|�������!w3*�O��Aչ�D;����[�3����#G�%fu���^��"�rA����ש�;ү�^��}���D^/MYvo�O�l�й�n��9if9��^�ſ�t��YP7�Qy|ڎ�VZ׎E6��㠻Jj�\j�`��J6Ze2���F
�x�N��-�	�·�>�\����Oa�eY|��B���N�]��J�Y��4�{C��h� ��d�A�e��v��O}՘�����A#O�D���w.s�o癚b�f^�/���9襀]�#�5g�@�H�h��d7��E}�/�DF�#}&Ks��񭭥+mE�w�Mؕ��`�O��rS����1�Ԥ{?���w˔Fl�%���#�i�e� ���Zl�����j�^'{��P2B <o
���@N�������É*��ᨈ�����J��Ph���[��"�Y�� �.ሥf��3¹��.����-rF)x.v���5���`e�?P���n�mdP�==�E��w �6�i��ʧl/���"#8LO�5��6�`E�7�0ۙ!d:�.��^�G#G���=Gq�~��e�
�X귳��R���ՊS�sf�4�,�iӍТ�΋Y�?������Urv:o�彍�l_xR�_l��}[Ͷ@h}[Co�8�̴<Re-ycd�����@�o��ܘ�m�l�M乁����R��)�6���ђ4����h�˶OTa��F9���8YD�H�����D�I����_��n�kn�ٴ�pu�W��xLV	}�Hƽr`����nRNH�ވݶ4�
��ָ���oF�'��L��:��{y��×�9��G�G�+X�'��FM ��x�8m�#T=C�6z�a�2^3�M��B�lXi:U_�#g�
���/�
��df���x�9N�LȂ��<yk�2-�˦b����e��G����M#L�ם�5�Ʀ^jl^�KF���F��ˬ�W�G�S���su7s�%^H��ձ�D�8�|��	��kؓK�XEl��]˚�G��+��	K����K������Zݴ��"Z�d��Ɛ���Ψ8���oF�X4z芭��ܐ��(9{Û�B�}��qw4l��&���4�5o���Η��V���9:��m�|*]$$~)�����s�N"��g��'����<q(���Л�BC�&��{�M����-���[Xې�G
"���)�^,�前 ����7k=�u]��oR^*ɋ쌽�,ΌQ��dc]��\,x���d�@�}W��|��;���Tr�=$�.�v����u�EW�c���AH�9�(,D��?ux��.`�>'��Ǭ����#��2���Q9�[0Z��R��I�?<��8"�cOhPO�6���~�'�s�ɉ��m����'|��Cb1h���'>7����:����?h��p�(���vhH&Y{C]ϟI���]���΀���lL8 �-h�&P�7�DG��5/yvh��Ж���r!@�f���2�mQî~l���M�8��ߌ!�	2�	*z�������|��l���/u�[�ts0vM�r ��"�&���@��ܼ4��d6_q�P��d�@��B.�F� N�D���ק���Q�ݍ�����; q>���V��k�(���1C�~aE�QQz��q�ۗq���۩Ω^49��sS�c��� 椠�j-�b��[o��ʴ�m��g�\���l�q�K,d�ta.ɷv��B�@z��i�B��>�]LD�W��cM a˻�h �"JW��z|q4�g�?uN��Q���T��*)c!M��s��X��>]�6�!���+��Q�5Bv$t��C�pn2�&.=���záMƃ9�W�k���M���_[�_ۼИc�?%e_CdYȀ���'g�>��y�<*��n�7S++����S9��T�%T�����dܕ�[Gp�&��C%��t��]�:�G�&!@��Cܪ �"�>t�d!W�dk�%_�ۃv=���0.2�a!ӠF���|#M0�<�Ĝt��$�K�n��2��|c�G[(�6�';�9�q�y5�,J�_�9�4y�`��!�&��A�3l��Vuz��:d�T���.c���͗�������+���'9�|Ӫ�����M{eeU�j>|8�4	��['�0���_����oƅ�V�&U����M��8��WcH��o�@��G����\ �7�n.��V
��|�NEF?FL^6��K��k�%	�H�(�
�;P��ܞ[0���e^D�)h����w����A�R�8����a��m�*���j��g}b�qϸi)A?گ����ţ_M0�������p�c髙�U:�����$lg���.MC��^D8���1�2Ѻ�I�f�]�UR�1[]YqG�I��u�%8��Y��Ռ��o͏�vƐ�1����tw0��
ht �_�����Ls<JV��u����ZM\�;B�a4�Rҁ!X7���T�<���I�����~� 7'U&T1�8��1�73��Sl��u�N�^�w%���kuUM��=v�K�yh�h�p��Ά��?��Mۄ����X:��n�6�[�156�ɕY�"|��Q88�U��$&il�rӷۢ�5��H*ሂ�F�Hnˑ��\�l����2��Tg�?3��K��ܚr*��LR��2G�*ߞntX(j�7�~�w��}\���X���-;Y������`��"c<tR�3�Wf��֢s�	V8��u��_��e��4��i@O`��&�]]:n�i���4W/z��\��</߸����R��(�߱�lx�T��j�aƢ	�~e�LȍO%���{u?u�I���]Ɩ�c������ߔ������ݜ��(C	'��uw��{��VÝ�q�ӞP��!=��oq�cP�zS�1�,9ǲ�\����f&���~ݞ	t�k9�FJ�0��b}�%�4#��:|�V���E1 UZ��>�k��MT�V��j�AR��g���i��|��P��5ť�z

,�WL���> 5�̗?�߬R�p�=��K:3}fxq ����Ú�.
&s���?�iS��6.�t�*J�=�p�������b�J0�ve���H N^�P�7�;
�K3��c
?��ȩ�2H������-���a�X��g��?w�͇���w��������(ݺ�;�l��53��r�����y����t�2�h�P�0_C���P8���L��*A6�/�f�F�T�Wo΀)u+1fp8NL\�V�G�9i) ����v\�v4�- ��W���0���(��d�*]"w����]Z�5���9��czR��-v�rwuj�C5S޼����1Y]v�rsz�d�����8(:�q���|��WJ1�7�:�T啿�[�{�o��44�,�� �#p�IFO�Q�E�dճ�r����<[��B��d�	�30$����d�X��zL�9n�;��N,��_wT�����=��ob��o>�Y��2_6�6�ڼm��BV܋ ��f��m�s�����'�pB��Z����3�@V'!�M�-ڝ@B�b�^����0��/@a/e-�:��X��M"���S�92U��*~dlQpd�{�:�0���ej���u�|�c	���A&B��FSUG�P9zl��a�`G^���@Y�
8�؃�!(�}r��3�&��I͍���zs5c6�ɦ3�������Z���g��Jq��P���y���2?�i���/C�k�+�K''�1G|U�FoLR@�s=MFE��9����Ӝ�q�)^6�@��.���C��-��3���-lq3���E"��<;���+F>��@���V\��Y��0����p��7�V�lj�qwz8��/��n�_��m�za���6 ��D�,17@���7��}|�k$�5��g'�o'(���YQV.�5y$,�l��bu�k�].�x�|Os�A�Q�K8����A��Ns�{�Kq ֦@P�t��4�d�����^�����r�Z��'�3�'ӏ�
<Q<��E1�i
W��E� ����3�����5�4����� ��� �
�g_�t(��3��f�m�����a�^��u����c�:�l�=��߽�k�x��w�pƓh�f����@��v撕:^2��q�!Ɛ��2��a!µ��yO"����W!)����'��s�Ut�����ț��g��0���;�|EA��Eoy��if��hq��3��tk�0�����1��u8�(wi�C -��<��c���A��Y z�0�#�cӍ3��>���t�L�F���?�:��U�Ze�,%\�Ԏ�͑.�H�~����f�??k>%���_��	��,���K��i�w���@��!e�Ќ{��J�_�������mRٰ��#���.
$��X����i�x����E�>�Ӿ��x�H�+����0����BR������
S�@�����'� O���+TQ��Ø8��T7�<&� YAmB���y�*�����������Ic�\ppc��r�'`�D=��Ӟ���y2���Ց��g48�����K�*�9ybA �+��b���/��!��<k�|�պ����&��%p�|϶�Y��w�j[6=O�\r^��]��#i
�+���O�ۡ���?Ì6b��d(S�i�..l���)���}4(��P`!31�H�c1��y�)\`DL�L�����LKUa�H��yC��3^��o�F������c�D7� `�����6�r6S��]n?8Q�P#��I;ľ$�/��:d�˗�UN+1�N����X�:Bg�v�����msV���O���m��v$�<a�>9�[����8�I� m���=��	DSV�]3P��9�uD�4�(�����Px4n���5��w~˯8KES���e�1��T��O�n�9�p����:RtS�@����w�i�w�7���Fv��� �u��|=N�ٿ�Ƀ�=j�E$)�7�8uw�&���e���q�)e�@,$��V�n��͓�!ǾM��G��t�F��\�pE���_���b��d9��uZ�0�>9��<�WX]�?�K�D{W��VW�v�Z�`����)�Nf�®��7�{��˜���{�3jp��5���`����z)I����T<�qf�
��w��|�mw�<Fk@�7, ��îl�O�6\8n%��d`Ny�j�� RT�P!�WR㻦�o����K8ȭ}�	��\�uS�_�����Gm���n&���T^K(`�l�c��_S������d6b��F�n�@F~R�50�vW��AB
ԍ���ۂq��ɷX�o���Ft�U�w"?�or�5��:��׷`~� �`��o��6��&I\�S�A�����0!����ݞ��0geh�pT��w@]qp�	��8�S�*�:��g����1�u����&�JH^<���_j	�ѣ\��_�	a���t_ ���"����n��L�ڊ�rB�� �É�3GB�%@3ϸ��8l�x�{��@�=��F��9�
9�b�����@�-�s5?�<J�c���!Q�f ��i�,�2�E��{k:Ku2扎2�m�/&OI�,u�2�n�!��
g��y�>n��π(�h��e��_0i���G!���uk��R���[����N�]�8T��緟�QA@"7��ư��'�{�\ެM3�X���B.]��%`��A�����Op'ջ��8{��\��h���Yao�t�aW����m��WYw����]	��%*���/\����f���`"��,�aY��,wnm�]:��g�ʷ��q1��΄AeF�o��|�:�pg>�t�[�3I����MX���ʓ�p�x��YS��kL��_�kPf�x�<3˜kKKe���y�8��:�P�n��|8X$=-8ʬL���*��A^����\�{�'p#�
��J%��Mse�v�����̰��I�Ɠ���F��ڪiH�Y������&���e�*�v�x�����l�D�q������/Y~xw�m����plv:sjz���$rx�����d�'�gLh�8pcǃ5���㔛}N.��q��q��a�fX|{�0���mt�a�H}�Ӵo�r�Y�r׎�����X�)]��8An4�D�����n�����⬫暟���Ȋ����W�4^�O\rLNV(9�#w��Lݾ$̣a�!��!��E����D�����Qh��4Ç�&�x�Vxsh��Y��e��/`Ws�"1��aNW�0 ̤0Ͷ���8�?	
�tq~9�VR11����r��>Y����m~-�I��<�z����_�k��{�k�Gpb\���'����c��?~LH�9 1'�55�IKTw7��F�z)��~�>������Ж�=�Ҿ���ny,Gf��[�(��n��_��� ��T�� ��&�+,�Y�,�c��j����r|3w��x>�j�������H��q ���Y�
��MA�7C���:::�Z9����޵WC p����`�[��i._(G�vG����7�wG�농�ĎJ��`����������l�2�*��zX,XXX\��GB�X˘Dv�EvE<�t�'���%;�b1��"��YFg$"N����ب��y���W���.yf��?������1O~��aֻ8yx���9HD�l���_�?sY�k��OlO�<Z��a�U[�>�SQCbbbҸ�Y�l��\�s��a۟��0�Gke��2��h�׏s����,s���@tΦD���z��z��E産�t���#.�E���� �,ݿ���p��X���W��,ⶐװJ�B�3�W6;;{|����m��C�~ZZZ�L�Rb��;l�滻���
�����o��X$+ݴv�\��މ��{����@�%赛�����}��j��ՀK�ǖ��Ѓ�q�9%�3o>g�U��L�Vϒ��mW��O��cH�6����ډ�u���.3	>w�j(^k���s���<����9����QV~Bbs`���#�}�i�����=$�Օ��ڹ#�� �v�~���v[s5hD�������x�l|���P�ӧO�۵B���������57?�'I�f(~�>\'H�cN����}$>ߢ����Nd9XT:E����5�c�:J�BW�<9�����م_SܹM��q�����FFI�/� ]�c�G�1��K�:����L����B��{bv�#ㄸ]�%t;� �P%㫳
^��a�p�m�2���s�Ή��^�vi��[���)T�epp$l>��r��+[��s�v���4+�1��V��1�M�iZ����pq����鮮.N��<�Ł��x�i��$���2>i������ ��q������f-�I��r�����M����Qt娌��~!4�}����Q���e�]��}����f�`be�H!遲���ߌ��S�m��_��.�ϑ��|�#;�K�l _��5�jY_e���E0,$Bx-��u��\q�=�Nl�?� x��B����l�������W�Y���I���JK�L�Go�n�VŴ�8��L�j#Fw�U]x�)I�ʭKG҄��u�t�^s�t�jhnRyy�����ɝ��U� ۟��L?#�h֑(�_bkHAI	�����:T]/23�,c��H�ɕ�B��V�'E�k����Xcz�'�����E�ۉ���=���4��E���9�����򠠠 �wT�uT����c��{'7�swvgN�:����Şb�K�9�;}ee�x��/_��k�F�a��8��e����s�CwX�a����������;��$���
��)�Άl��aέ�pt4n���:%z���|�U]N��w��גۨ��Qv\��2i1T�G�Vjw����r��yb�JɁ�^T��XM^ja!w4�����Z�G}>R80dt�&�ݭP���N����:�X@Spc��$^w����ӘGz��c���b�Gph�L��t��;�[$���>fN}-�ăik�ͺ��"P[w�W��d���`�F���i�i��V4�o��w��� TMMM�~�V,������3��X�rkR�vW�s'ܫt��/��Y�*�Tnh
	�q�TQ:�����P�3�מp�Q�$AC�[%�#bâ]4�9'bm|�
�UH�Whis��(y,��RN��3�Y�J'�طq���=������f^�dp��Dm�HjU�����#�$�@T|Z���y,�og"x�#�ӡwd��k��}����)�I�EN3@m����̜��Z�[�/)�J����q�,��Xa{��
������ҍ^���M�/ȧd�w��v�����x�������Nw�p�]� �f^��Ǻp[y�C�xl�p�OTtql��A�����b8S���K�z��K��|��#���i�����^�X$	��+���A�ߝ'Hм���W��{+�*���1�^<�\�(�Ъ���a^�͏_���=37	������Y��OB��嵫P�*����h�x
Ҽ<�d�^��^}V��ӷ�A8,22R�e�d���|d�j��aܵ�h~nnu%�Kp5�)?��@IQ�,>�`d��9��}�.��8�� �e	/�S6����ݳ7<h]-D���@^W��sqA���m�°T�r�m�855U�Ό|;7�!��ڦ�p;�ջ�pE?�ԋs@ڴ@v��,�e��i4Fܚ�^��Z�k��՘M"�R�hUnߣ��c���g|$獭���������|t�x�t	��t�*�M��]�5�����i����*~Gǔog��g�d�EM̱g�  �v�ݪ���ٌ�ʍhW{Bυ���GUl)���@���/|�'�ːe���:^�����o��c`b0�LCƦ��@�@����c��cB�5v\k�H\����$e��M-Q�J=��	=u�p��"k�"ʍ�G������4O�����5у�lJ�c�v�m�f܎�݁�m�#���uWt{� ��������s271���pb)))`b������R� ��M9��W&���������l8>�b� "�@��M��n�6�&�]Kb�`l�N�oۄ1�Ekȍ�^����C���"�Q��^��Ғ��i�X��n`�b/t��0o�R��?n&Ђ��Н�{�_@2�Jr#���ݷo��|�������ɵ_nɄ����g�Of=��S��˴X1�U�ck�C�Q1\�<e�_;���^�5F��>*?;/�$��Jl�]-[+.�Yj�������{���+TO_&xƈ�~i��0�b�YdMdz.3��F��q����} X~G�)�'Lt "�bW��E��ҟ�P�&wpp0���]���-��%�����hN ]N�A^Hv[�ܩ�z�P��h�%@�����OT��+�BE��2_�a���(Q*Q;��;a�I�`���v;O.�gR�kC�x#�2Q���K�~2*�5����^r�Z,���;p��D�8u���� �M��>O������z#̵���� ��T��.�%�����>�G�5\`G}�.��"���[��0d��3k�1������,�\C��r4V3++V�'����h����I,_�\�0�����Z�ͬ��_	�Fjt���SJ��O�=L�X����_V�]Y��%���EO�aǞ6Ԛ�ǣ�\*s�d,�����f)��-��×h�,@L�ХE/�#����8;��uP�$Q�-�Fq�lnZ��������W���RT����B�MC��6�**I�?��ZXV0K^"���<;Q�(y�fS�i�Z}�D*�ʠhyJ��?|���B�
������ ��E/!iH��N=����)��^R�T��,;�H9Ȝ�i�_C��{���J��f�����#���'����Tם��!ͤ�a��C1ϝ��;{=�7\�PX@��}w�~��z�xd��c���n���.�k|�sKH�V�%�p�@LM
|OZ��Q~	`��0m��լ�87V�|5���t"�;���G��R{Ǡ��oH��	��եu��l5�J�bn�M�1��2ۘ�w?�J��ݏ�>�0�Q�^�%�w��X���ݷ�0�?���1**J�43�
.lU�XӦSl�c���-�SAج�m4�}¨�f	a�HN����|��Fc* ��|�.A()+�XJg3����Ks��7UZ�m�.b��2?���:����XXX�;��q^9E�.v��ʣ
`���!Lllȝ+벧Qt�S����#w7����?�@]��z�'���B?��=�!��,!�	>Mש����齈�(c_<����
E��ýG�n^�_hXzCt�������̷�8q��1b�Dי�'����?X�[����a���=�m7V���N�C�rss��p��B';i�G�Z�Q�L���U��^_�cV �|ϸ]C��wj�v��G�H�!�7Vr�F�E�G��5��]����7�E(�{��� �Σӟ�n�� ��8����yN��W�V��������k��)�l*�ţ��eL��=d�4,������N6�D��\�ӈ���u ��ƭ�̈O�?��ၭ-��k��jzs�\�Ǻ���M��-���6��k� `�.0T��s:z���@IQO�&44�7~�7�1��V��j�m��K�z����oݻ�i��r{o@�d O���^V{��}(&L�{3�x����G���� �6�*A���i��
�19Q<�ZC^�p�(S�ۂ��n-������|��R�f<�!A+'p��^�o�:���[@��=-v�h��u�H��F�&U��T=�N̽����,��4�IwI�d�
�^426��2�.�Z6i;=7^咽DM�Z�T2�dk�px�'�@�'�YK��T�"��5�˝,׮�:������D��
��?ϰ4#uNk�N�Dο~%�W'�P_�f0~4������P�Q�v"ĥK����}����� ���ڵ������#qmƤB�A������r��^�y?mP��*XU5S��?�P[y0� ���t�IL��9o<o��M�%��HP}c
5,���2��x:v����%P4��1���˯�Q�^;k/���3¿Vп�I���73=]��m~!�D�&�΢Jo�_�	sΉ4/�?ox"��^⍯P�jj �b#9^�X�v�JW��_��xK�s�am�K_)ƗS��^�w�L����֯m���[*2mbV�����p0�'(�~d�W��\�$�uШ�1~.P�}��ff�߳�S L��@X�_C�5�<�W\F�)?��������D[o)y��|'u4������n�k�*��(���c�ySʢjq�q�9�yl��ĳ�mU����/���hc�Ƿ݇�`ܢ$��^`����1qG�kׅo�^�E�h��@>�d�z��ݨ}���J�j����wr�<�>�#QMYlݫ�f�_��vR��.+�6yE�u2�25��I-Z�5���y������'�����u_��%W�]�N�,<���C�3���s��|k'��O�A;��+;���������μ�2�Z|uƫ��+z���8�`�����3{=�� �I8�a�[�>^ڎ8O���M����2�`R/�����9�I�HY�n1�\*@���vuZ�L(�E$:�`�x%�W�GS~/v�͜ ^vm�h��ƍ:)��L�\��O�[_��
L�}p�Yi���C0���
��k�ɧ�D-z�u:]���L��O
.�,����>���������8��(m���k ��1=}hBK�ӎY7o��f!�.[i��)�A������rt)���}�|����h nc��Y>|�]#{�x]o_�n����~� ���v�-x&�D���gԸJ�oϩ4y�as����N���ɠr�L����e�/=͎�	�oDv���ّ��k?��܇�5]�=
k�l	�Q�XX��]+�+�F����yȁ;����Н'�>LT遏(�0��TJ8aH���9� JBC��Q?���b{��+[�-�š���d[^5�f�s�?����b��9�܁#]���!On���nwǻ��9l����,o�.�>}w0��_���Ł��n5�C��ybv����,��F7���=<�9��}�뺝H�A�N���`4Uuu�jO̅�j㶨Ɓq��1�e�� Z�`F�}�Ҿ?lU���~w����'=f>w��2��x2�D�����B��
�l�m���#/|�O�w*�'!Ѳ�zd�6��J����o&��-���@#s�
�C{�n'�@N��S���i-�L���ȵ�M��}
��׼���(ľ��,��0�{���0 "�UD�D��̳dH�NTm[y�� Һ}$@�C�KG
'����n���i�.R`��`_R�zXM����8��������"�b|q��ദ��4� s����F�ڨ���A�mN7v�E����K�&J��ag侴�ueF���O�	Td^?�����/���>\���q��>�p�h���.�'�9=�����Q�omĖDN�֘�s1�8��P�J}r�s�v�����I�������L�c�����u�W�.iXy�1�+��M�0�Z5����c9�R�54�<e~�β�;�Ґ%�	W~zg��7�(�.Um���^l@lQ�8��'�t����/>���r_�~��Dӻ֛�V�͸7�i:����ً�2�ʦ�5��z���;�[e��,�U<��l#Ǘ�&j�E���Vz�R�1�Z�E�ͺH�q�}�b��p���T��'Hh��R������1�L����/~2S-[�A����ݽ�Nse��Q���+�'�6�^'(���з	xu�����9ר����n����F�'��T�i)Ǹ�	)ȩJ��!�޶��ab]eǭk>�`ڕ"njj:��g� ٽ7����<O�(�z��j�������>��HO2��7M�s,���,�	�I�}@��!�SIW��p�.�
M�q&b�nFù������&���~w��5l���)��`�c�M�S�o|��ds�R��u�~��	g]\��p���x����gU����J}��������	)lT���Ue��8HH�ֹ�X�W�������������}�N�6J_h���5�Ƶ�[�N��� tz�պ���PUU��ifn>�(�#E�\�'{BԹ���yG�~̫c��%�����С�4�O����2���$K�j�U�b�:$j���;�c-z����4�`qp�l�ݘ���ǾbR�>\��6H::;wV�455u\g�W���&��)���:�₯�A�!�OF#r��-܈\9��Rɬ��?ʾ:*��^P�c�@@�[���F��.��N��N�.�����;���{���}�}k�Z��{���~���9'����[>��K��R�
�7�R�{ɚ��pW�=�7kV����pe�����O1a4��yD"x�xY�ևih�'��b���-�C��� �Z���)��+~<9������N��6�c���3�o(���..��8�<.�诏9���j��?��H2�SST1;_b@E������y4���v�U��M=�QV��!�F1����V�����t\���=I�����(.�r�4���]���xiw�螟�%W��gH�?�~�;��ˉ#l���bY��H��
fm�=���t�~�X-������x�+Im����|�}�A���I36�F�y�`��
�J�Vܝ?�Չ$���yH�Eu�Ҁ��|����Z
>ĥ�	����Ӆ�#3��^�X�K�D�,!���WFqo�}zi�8^f���{��!L�Aco{F#��6@���=����a�DFu��m�n�9��XT�R�k����dE��?�D��<�T��X�=~���� �&>�r��L ��JB ������l*�8���]��~��Dk"~g[���w��8Ƚ�E�:�l��5~��68�#���C 9��䫴4㔯I��w~x�S�y�zF`o~i,���	}���	����'2f����}�py��΢#0�|��9r�맃0�x�]����(�s��)T�������
T@�{T�k�G���=�⧮�	�1�L��~��F���bki���s�����;ӹ�;--������y�MU�&&�N��K>�/�ͼF��`��bP]z�),n��1˦3�PL��������X����v��g�$ɝ ���K�v�oo+LQ��>�6����D>;��Q�W5��O�����Q���.C<N�%uKf�YG��I9l�_P�ݻ���Pb2�ǵU���NwjoW僕���nr�+V�{r
�b����q,��c�aRo\�_i�}�=IR��}򾡥�ݘ����e�ͳ�p�zʩP��׽t
�N�C��b~?11��q�tņ�Av�����D��`������I�f	n��B���(����49�!�����[���mQ�]ulz[iAH��s����mx�rh��h��Iw�U�9�0{8s�됖�n���X$|>��р׻�i�����V���$�-�h-w����lt78�B�	��{߳�qG�,BED;:��s��.P���߬��G����D��ݵ�v�s.\�GMș/D��azq!����-�ta�k��"�2�t��q�*/gs����yo8�Ӂ�Ũ$M��}'A\0��A�U��[�gjͱ��������oÁ빧_V󢃼ff6'�����U�ƣ��K�h�J۶��`d;��@v�1��q!b�h����xY��d1��;�y�[ M*�������x��L�8�2�GR�䎳�cx,���(���h���/u�� Y���H�k?a^U�� ]8Z	��Z�H��v��3�ǭ�
,��6�+�	.��dt:[%i��\�l=is �_��8:�32��V'�XQ���ӤN�tq7���sK����ċ�ۉ#@^^\d�w��A�?:qվo�256�+��h<^�'��<� ���ZA@z߸��0�v�a���b�Ӡ�[c���H
.HD��7��c��GաҜSxP
���L�/o���ޕ�����q����>ɼGR�ᴴ��U���/ͺ�OU&i��oog�cIR������[]����� ��������/�y���P�8���Rd�[��uk�?eg���a���h� +ڍ�	vW������ގ�9��d�β��fh�ֹ�]y�a�J<V���A'̩N	� )5�v��ao��ս�*u)A/\��5~�-�0(\?}�j�ύ�����P!7KH���4 �r��tooo��o���;K�� e D���?��B,�kd?g�ڈ�ѽ��-�+����Se�ZtKw�<��/��������@�@�մ�J;@N�/�Q��S��h��MCAR�l�  �*���9]�l�\��LCI�*􊖖�_�~�9�hۤ����]�6PN�Q��A�%����IR���g��x2	���X��/I���d���A�
呪�ת�P��(��
Y��~�ID>d��x����I$+I.x��*-��� z�U\��B-<;�������x1<���A$�@�)IŲ>�;E[��7U��G��΋qg�ʇ�\�*�����/��:���n����۪�s�9��X`Tm=�3db;EZ����hMSX�4/:�h�F5�J�Q5#� �_����^^���"��3C��*�8�SR��A[�1�k�Ӎ.-���CU�,$<[Kz~�s��Pr��&��sV��;5.�z��JG�uwu�7l�Y�^�����\O(o����hD'�P�Hb8Vl'm�b�m�<}��Ư�;/�ʜ(�k<PH��6Z璻z���7JN���?
X�O#��{��~���.�~����\�����oGNm�s"�B��8��Hnt0�R�gV�6�-�vB�����-�̫�8..��E�X��p�`����Fn �w�ޞ�KPq� /���E�����}�ţǫ�{�A��z�K�ޢ������C���80���8^����7� �8b�N�+e>�ď@�f��XB�GEK%�����`����C��W��k�o�6?M/j�]�ԡO)O��hL���t�R�����x�P�w��l�P�	�?!h��'���y;�LMM,=N&�?�3-��7���.mD�W�N��3$��Ƌ�{���p���j�-^R\�<�EY�|�6YM���eGǷ�l8�����D/P�LD����a5�<	��>�M�U���L-�D�n^�Ի�ܼ���A����

�y��{�K`�H�8`�L�3|j�C��K"V:��Ǿz���Z"ל��h����6Y+-eVF9+�üb�b����}����B���Zi�.�HIK�ԗ���f@�숞���5��a�j\?Z��ɩ׀��0pXo�s���[A�R�m�D��?��ҁ�K��3��Ӑi�T���'X�PQm�O�NW���(���pX�uGP�	U�;�#yJV;��Ў ҡ� ����Gs3@zy�� ���o���v�M&"2�� ;=�](�	����B��9��A�V���Ư����68*W\<�[u]|�Z��n���l�>$"��7ع>N%�8�X?����{�S]��;��w�;i�a_�FY8���ZYI�U{��/�OlxvA���Y����E�.�>�Sæ��X����A��M"�a��o&V���7	p����!��}j(T��ߞZ��K5��:k͡�\~���7
-8Q�d%���& �P�r!���K��O�����#;Dl�6��M�#!TƐ
�/�K��3 ��h{�f��v莟wq��<�t/t�D���l�����1c+��e)t��4L�>xLr �n�t4����:�.aY�oG�7�\��<���o�_�nOO�߄.������d����-	C5`�a����4��j$jΦ{�g	��*0�;e�yI=�BTH�wf�����޵�s l��Q�
�׾(8K�σ�S�$y�t�ϭAx���d����a�'ՠ'Q~\}����ka��~%zЎ6?ܡ���#.�$��g �@|2RE���#p�lY>d���[Ծȶ	�1X�r��W�ջ ȨC�[$S���;�SSfn�*xP�Pd� �|»"l�NAϫ��O��+����Tb�dS^��<,����~�=�à��à�@�[ݻ��?#{X�FU�s+���>����o��/�vi8L�c�2� 4���U�9jcT��&�Í&'�@u]�!ujE;(p���FaU��8���X�6 �k��C7�b5/�-&!7�~S�"l�����\#��7k�B����I���5�0ĩ�d>#����3-�dL���1�S<|�r�V�ͳt,��b~f�FM{غ�Vp1!���`W���7��Bg���w���R����-��x{L��/���`���fš]�5�k%�&���ˠ/)qh\�}�� �VCҜ�)���X �4	ؕ�}�޺�X;��T����_�ᯉ�����H�M��e��P���Ο4i>�ᨺj�	���s-��̓zL2.fW|Ff��˶���8��|g��A`M�� S^q�FY/ݥ���^�Y	�>���L+��%O���w�	�4v۾xsF����َ��HZh��6����A9h��?����w�P+���3�z�"����ݵA 9Z �E��p&�Q���f���#�u�j9�!��+����A��ܫ��<���� ��q~

$ҁ7E�l��%��fCn���A�̰/ �L%Ǡ,)�)�4��i���MH ����9�V_�\�x�9���. %8ںpa?��R�2�n�2�&p������g  ��x��I�� ���"w"֏�O]�Z��U�< �uJI�VN#B�8v�����������d5X"QTV�w�Lp�@'i�)�[�>|��`>cuh����ŵ��#'7�o𓗃�� |5)O��Ld�d�2 �/�Qs8� P�@P�d�p��a`�g����j��>I��^��W�.l���KYi�V�p���ǧ����b��$IMyz}a^^ޘ���h�hQ9�~��71��i��~oޘ��x�	,�������
�^����1B%=�4��'s6F�b�\� �bl���� ���>z�0�2LϐP9�1�-�Hb��P`<�;���,�w�Kp3P$ƅZM_��+#��,�^�������`D�t9�N��N:���������{��%6��N�d�&���AsXjt[�rԌ�&A�n�C����r�U80��F+� �q��猫�W«�'��J���B��[ �{���@Lu��������"�	���b��t��	����T�d%E�6 ���O_V��>M��7| c c�O��
2w���}��@�����jO������T�~!�Fc�U���kEܘ-��@�	ďd5��q�� 0��� ��>1qI��N�	���4��@e��V��%���``c\�������#���'88%;�@�AK���#�n4���.���f�~�����\:�5��iL�ڕ���I�
�������-�������Z���A	�f��V�'啛����� ��3S�~Aq 7-���~ e0H���5���*V�6ߣ��2��t�L��$�A���Rf�ƹH�O�nG&oe+-��'wf�:����{�.��)Y~�b�݃��>'k��������5����QLZIeN�*��Ta ���^n$���ട������Ӄ��i�M�u�њ��3�@���X�٧� � \��\�9�m �p��yW:M� �G�V+keƒB��[��J�^k��s����bj�Q��py%���i���gacի��POE��̠������r6�n���6�n���i:-E1�`왿me�	@�����	�\�� �*�i��o��,bV�$�ܩ��~�k�p����aF��L#��@���E��@n����T���`#���ģ��,�Z;L�O`@0�Ouڷ:㧛���
X�fq�_�R�Lu����dHQ a%=-�i�M�l29��'a�]��$gZr��P2�VZZ������>.* ?:s�N C�/h��ZM��8�Ef7,�������z�(�Q&d�c:��I�x�j�(Ꞿ�w�
�mh�����1��C��7�/4O����R����.�&&�wM��e
\g}�%6�CT��`"fm�^C-�����ۊ�K)X�yo���A�8k�� �8�E�PHKo%�ؒ~���&�f��� 0��Ɠ-�"%��dff� ��IDʡ��zzz �Z��tһ0Ǚծ1��1���D��s�{��-d.I�8 ;�_	��w��\m�x<�79waV�Ţ�H�ck�k��0e*���4-� ��h��tHC���U�hύ1Ў��, �C���#h�5�����``���w!Ц:k�̑��(��޼�,`���2."�?�� ��,z�U��N�R�Q�<��د=?^�sv�6�e�uRR�U<9�Q��ičLO��h:���~������߆�Z�����"�}��KQ�����2���@Е�}�C�@cjb��##ZM���z����c��y=��T6%j�E�Π�b��������gq�%���������{Xb�6ȵ��>f\O��� �`�Ӯ����z>�4�W��"��ȱ������ı�=C�k�߱/�	�".�SKJXz��AV�\�Bg����e��ӫW�#|c��� ���b'�>N��c�D�'|���B����G�GV$��#�b&�	����+�Ʃ�K��C2777�����ܘ����_癞ӆ��#��	SFGG����D^N%h���ʅ�6���E5�q4��2�2& �hj5`j�q:�4�r�������������(({41K���M��k<CXRs4�~pAT��q��nC[�������ʅ��#�� �����+Eīz���9���w�3 �ϣB:���H@�H@�9`3Tޘ�;�6�ZL��Ow�%�܇ ��a����M����M=��7�����x4��D���2����J������B$©D޿�z��5�uq����_��e�c@���t���D�dL$�J�����cs��?�@@�f���E�g8e��| �Է�
�̮�Mޠa���Ke�|���X	ҋ��	������Lǒ����?~��L�l���`S�V�QL̘sJ�d���t�� ���$���y	]Z��� ����y�Y�[hӠ0�Y]�����6��y��_	&ڽo�^��y�_ɩ��KF)������<����+��JE����L4����c���<�F���{n]�iJ����;�ED�8�i��Ñ(A � �W.�=0��\����s�Ü�ZI���FD��g}��Z6�j���|�]!�q��&~5����SDX�c��\��~��b���8'�Z���J������7��A:�%�c��[�yJq�,��&�M�5�G�3 ��S�r=���9E4��
�l���C��8����j=i��s�o:���1L]���V;l�wgA.ic
�zy=e@]{��c�)s!�H�L��m��������μ�(����W���&��_��=��ޘ�!�ٮ�ɯ�H��S������{2�m^�Zɋ꥖H�OS����3ӬE�������	��{GdA�"�7Ƞ�F��F��?�f/�x���_~���;*-�X�|Ҫ7s�'�{��f����z�Fڷ�N��TС��][F��a��~��Y�`���]/{�`�A�?/��0�~LmaڵBW(���k�����UeX۸�N�c:��p���2�^.�ذy)p�pnu����v�WO����o�]8��x� �⨴}#� F_d����,^�b��g��q��l���P!u|�z�b�!��~͞�W�o�����l�,��'RS i�߼SX�O*�\�&Y�ޮp�t���q𒔔�O��(�%O�i�<�5֐�����h[�7��1@�y��((��-=a��bŦ��խ'.m,cM`8�'\�+�/bu�`j�ze�UW�]H1M��%���ȃ������U΅���"��'�1����#��6�ye}!)�^Z�������â��A���i�����p��X�W[J�OM���	��f��]D��yV�|�T�����(�!�镞�9k�T�ǴRri�џ6�Qp�����W	(fm: �K�1|�W�7yRn��.�K�8u�<L/3]:p�$Y�i��T�`0O���B�%ý�k`̣��t�[�1����~b\�����m�jU	�j���̔O�;��&`f
���ꁁ9�Z+.�ԟ!;4���?!8�#�@�A�(�}/�j�r������Ɯ�,d�=Q�@�?6v�6�*�&+\�.Y}����k�Zί����8'fL�1l9C�N앶m��L��Z�]V< ��v���.����oRT��	V�dVm8@�Z��0��hȧ�
�R���I�=݇Z��9�Loy�_���OFd���[K`6:|ۏd��^��cvb#�w�5�*&2z��_����
.�#�'�@	g�P�Ӱ�|���ڪ,�spL�G����u�����6%���j��<e���B	GN��VdZM��;%����'�޶�d"��ģ����\��LPKr��5P4]���=��w;��Y�]럏��@rWj͋�OS*���O5g��m�_v�+���'��eny�AA� �,N�`=��Q6e������r8HSꏒb�7�oWh5�s��z���1[��+������Qҥ���|��+�}lB�p��z�����(!\�˖D�[ה��f/�
T�z��f=#�Z��j�pq�,D4(��p5ڼ�t���|��L	|!n'8���r>?�����A5��F�6���ťK�b<�ItG��A�j�����Rp�&����S��ت28u:6��J�
�[���<�mL���*j9�@D�:��po��2 ^��3b��� ��L<��;ӛ��/����4�L��)�k��k���!y�*���%�ɑ����^z��
W�Tᵏ�!um���w�8�jkK�cL*Ρ��*t��C����ccw��K�G�#c��/�>K	&�g��Cv���j�?�-��N:������tmv��zh��i����f��\��~~�qj�ᙦ}E�܁�ɏIA�_�8|��(�X�qk��N�+�f�P�yY���i<r�.�����&�o<}]����G� _�������Z�0��D"�>҄%��-�
&˭2��2��UE�"I�v��*T�D�\�h@�ݙ�JSuK��:�y����"����'P��7�M�iɤc"*wp�9�@{�~�mf�c��3N�Ze6��𯯇��<�1*ac�c~J�Sux{��kNzMԹfa\Y�	����ڏ�Q>��_�B�Aʹ�����5"��t,#6oS�CS_>sJ�9R	����	�%�k��=!�M�о��N�޴�:�nrr��V:�E5�!��1��7v��k��H���d)&�o39ݞ3z-�&R�Ѩ&�S�TBH�>�����V���mI��䍈��{�3���b7�8�uϔ�����F�sCmE�������ő�-��L!��Qb���#R7��C��&5nx��v��Z�â��kr�a"�`ơ��OFm���B�h��k�_�&�6�����~��r;�m����W\?���0��xም��i��Ӓo��ɍ���IS��i!�*���PV~R�JܕE{��M�:�O�#r�t��3a(�l�C��w�Z�>,`���`�gs�w[�������\����=���L4T�l<��b�������w&����1��:��qf�ЙC�xgfz������GG��%s�=�Vp���]����ckWW�t���o�Ml�+���>��(��m����b�j-o�+"|�QhF���/D91�=�1��VO���5M�{���{YH3�&\	!�����`���q��\���9��8; ��^���p؞H��j�;Zv��n�����.��Aa{�1�q�SF�m����c�Z�Oڠ�]3���U��>��p�ٝ�ug�ȪF�[�!�= � 9��PX^2}�%����D"���tul�����B�owKn�(�-���6H���9P��P�M��Xu�`l��7��凮�6�`*��g=�V��*��ay�ݎ��YR]�`ƫc��{�4?!���7��IxB���!��WC�mP�7-��f󿧕���9�KI,��j�u�L�
~�v��n��:��d�u 	��+�h}�?y�qg�__G�FѾ�@Ӫ���2��l_���2s�VbŎő�������$���ݽ�����&�����=�Z�c�o3�ZH�?JG�/0�?Xxb=''2z�wnsk��]���@�it��,�η��RWo�\2n��vq2�"ԌY�	�x�4u��ac@�b���[֝�AN��|���zn0F�S�V��+G�Z	l���˅I��17�R���e�勳�tH�{E��#b��8Α�*�����B�U�|u�h+����w~���������mGN0U�~����.��ʔ�2�7`�CY�$DD��ɵ�����n��G{ү��$��>3�N^�e'}/����p���wo�7��7�·^�-N �p%SAWڭ��俖�)�trσiyhЩ������{���k� ��>s%����?"0��Ƃ������G�i{�gv̇}�59����6tm��)ũ��:�m�pw�'_-�Xߕ9AF�]���5�מ�N���|}t�]�F��u2�}��*����<��0n'J@�ȉ��5gJWe�~ܨ	jH�<2®�����/�:�i7���x��m;�p}�	�U��E��|�ؒ󀑢Ì[�V�c�R��*��
u����2�~b��*�m�qQ��Q߉̚�l�`l���&�2���+�?-�1�/,�"���.Zo8���4?	=�����&�K�J<(ެ�xH��-�G�nc&:���Zؚ��Y��99���e���]�ځ=Cv0�� �Z#�"��m�mx�4���K0~��8i�S��>[*aO�JmH�;�}]5�ӌ�E�nHL��0��<�F�W]�9��z����!2⏱���s��JXH*�ۇ<	��Is6Woj��-�q�8��R�R�Ȗ���21q��#ǖ�����c˻����XXV��ٮ�����;��XN��$�͚;�-��U��X�Ol�-��<�2��3m�Fa.i-�3��^h�xO��K����z�/~����35gǖ!v�fqJs#��4��^�<r�Oj���o��
�ƍ�&Z�~X4�+�N�u���z@���K���N<9���\�?"k�38d%Mv��U���T�bg.��m��W������9âmE"e[lƢ�):�IX,;�g����d�Y-uy��V+WV��W6n{��8��:U+,,�E��W�m(wߙM���x����{RpR쳪p�p�Wr^6�lH\1�g�fƲ	9i��0��g|�fłԕ�g��?�r�U����@lǂ(��W˓�b�{[���C�1��W��Xj�D��Y���d36�Z��ڪ�3�Q�\�3s0D~n$3�v�>�QQ����怊,r�*=��q��]i�$%��k�)}6+�B'�#�PV<>��|��-ru�Yr�7�b�����n5�F-ֈ>���*�����V��F��m�GT���>����~���� �w��#r�r�k���^<g?N�D9�ؙ� G)����C\0��ؖ6���ki��fbFk�M*���D��8=}���Bn����՝V�H}6�P���,jרD����h�~���gu-�LE��%������08ߙ�Ht�k��M��=���HyIٱ� ��RHrH�[ t� �k����;���4խd�U��Aҟ,ז���b��G|�z�n/oߎ)xFJ-�r"B�O�3fe�:-vp|;Nd �8CIDk�k�k/2\�vb%��n00֘�+6D<�$�9��%�b���Dn�7��8T3��Σ�9��x������+���QO�O
�,�]xT;��+�a�]����ϵ���tC���!��8B$�����2#��o���,��lI]��0���Nn�dpj�F�R��(�O���ď�{���)>]���S۰�J���f_��,-���T����3���[�G	�� 7�^���v~��X�"4�,k�������`��@eT���M�#'.<?���k��N�oZ ���G.��1�b� ��j�c5�L
�v�o�Ww4�1W�#�5<���Yk�8������,��d�E������V�]�#g�e_Ѫ~�rti:�*�aT~Z�:Ms�|��`cb�`�h���}�������Ǉ$�O��B��S��uV-^�M~[ؠc�'����3[�l���;��	ɋ�vad���u?�-kb��S�jq�~[T����� ���4�p8-Y㖐��;���.@�ɲ��RT�t�\���/���4,�@�����]���D�%Q�^X�S�|w�E�����)�����EJD������^��}��|�!��Isz3G�W'����
�V�^T	�+��J߄��{bb!���y�3�@�$����������c�`���A�x��!���8��Ǩ�ݲV�&0��3Sɛ��&ngJK�Ԁw,��8�V�?����*F�X�����-ڗ>��U%t������9�k
M��n��Ԣ���c�L�D�ˢz���ɷ�|\��6\�� �Ӵ�zMǵ��7
y������GJR]�hu"����#o��!ڮ"���Jr�`K�K�"v��[��>��2޻���]�z���"�kL4�}�L���=�?I6�$�d%���
O~\�*@�"jc}������*6`4�c�����T��nV�

z��L �l���=�1�]�oHw����ɴ�e^z�s�A�����O�Ղ��P����+?c�E����.�Τ�����xS{��+�d1�����VU���s����0N��ه��j I��|�:T�ῑ�]+^l�����A�Rc���pt1�I�2�
T�|�wG��ihl�T�`���%e	����߿���Z:Y�?׎��uo7��d4���(�#�Vw��U��J�ER���0|�'�� �D�Eܼ�*��#�:in%|�tz���}r��
,���Z\"�w���v|���i�9=�{Sx�:�`8���{��99iZ=��b�^�L�x�p�&�����O&m�^�p�2�S'���D�[��,]� r��{�Y�XՔ]]�@�0�_�h��L�q��x�!���)�K��h�zݙ��
�������g s�Tnx�X��ײE0��|����/������������݊�V����P�HHe0Cy��x�	!�yٜu/c�r���%��ok��v�������r��ߵ��;*�o�6��U�5y�J�xR5q4���훨����Q�f�p��4����u�0�G �5k�7�(��EC]��)K)�d_�n�kB�y�ɤW�����Q?!���E��шOg����D�\���ŷ2��t��h{��80;Ns;�%�uޟ�}@t���R1�a�˨��r�t�̨[�bw������ok��Ω��U��1�t%��������:|*�BgC����O��n�<���v�<�I
����i� �1Wj [	5�a���O4�*|c��~�b�~~�ls���~�E��k�?rTK�l�3c����h���Z �U"$�8�lh�0j#K���т�}�B�a_Ử�#�1�ʽ�t&]��c�=��f��@A�&ڳ�۠�kG�m�B\ă�7�]�Tζ-�V�t!��O��t��f��`#��j��t��׽���(	���	z%�w!�3�����*86�Zit��f#q�ڕ�`�ė�y*3�����c������E����L���e��ʠC6���n��g�Ќ�l�������*ԝ�u=ph춬�u-�<MX�E��%�@�:h]7��F�f5[�s����ʢZ���o:|���z�%w���n446x���p��$*Sa08��To��k��4� �N�34��墪s�g�Oq]nt��,\4�����޳�C~;/O�T9߶(,�f���̤.�?�̠����Ĭm0%$e���42������;����\	�1&����I�D�	���*�Q�ho֜��{�D�$�N~p۞��_}�ϟ�r�q�W���uLME[�4�W6y�n�nt������� .���FOoE@�}/�EϬD��XҕD�O��\���]���uѝ��* �������B�ۛ6��>l���^���߁ ��C���a��Ʈ��*`)'�n��(��zOOC:W��ȵ�@	s��#}R?B�����jphJ�[��ivDN)M�0;lsg#���TR���sI�Ñ��k�miut)~W���чs~���	�4<˼������������[=P����A��I���ŏ�x��Dr�( 8�^%�,�{�TS��*�f:�${\�&�G��pI�ǕA�^Rz�Ŗq'ͤ\S��Z1A�j�ϩչ7�4^&�د�6q��l#��
�����U��G�[�t���5vr%���X�ǽi� a�y)ۃ�-�����??�v�����k��r�tw����?۴QB�H<����p(��,�]��ۮ��xrQq���1Ǔ��d���".�r1��^O� ��C�|v�IQ�q��&�Rc�'����^b3��?
��c�N&ȫ���¤�8�h Ⱥ���nC+~�A��Y{�ͳ���GvtnZ��5O�<��3�U��u�N�+= �� �*l��{.�e�l~��o�_��1�
	�]�1wv>P��Q7�x���� �Ѳ��(��!�S�f���.b������aċ�v���G�q����G�Y�� B��V�������6�'l��B.���}y�f�<)3�(6�Y'�����7!�U0k�F�v����Zd_	�����>�*b�y�����#i(�<Z�kY}�v$�!�;��CS��z��P��2��4}y��C����
�ے��,F20��Շ�^�<޷��)OH���'�������=kd�#Q1�}<J֬�>']��V��
7��xò�v+�,?�,9��?9G����)��)ү����s�,t"ˣ�5��T��w���iڵ�M�&��b2p�/���1?�A�/�����������l ]q�_|��*��N�C@��A�Sp8C�)�6�nx���oʆ�\���V�,|G��s_�(�j9d�`�_��=���n⇝��D@��k�D�s�d��i�����ݶs<^�Gϐ��|1S��t)�O�Oǅ��0w#�׸�s��Qd���v������A����c�?{����EThN�chm��3h���_��\E�Ҋ���7bցN~��������Y����(�8Q>�`͉QK�@�hw�����	�ӝ�O�M�OQ����i#����"�r����,������_�L�e����L�FaVAf��ʛ���0�&�]���f�G�v6�c�jզ����	ў� ��{�T�g�����Y�Ky!_B������z�z��w����`�ǝ��ć����
͜����,J�'��ǳ38.6}-3)vWd�Y��Yb�6��Vd�!Z����Op�9l��������m��/��o&�_��S��#���]���d�w��+���� mܟ�r��ȼv�����RUN�6ۈ��8�'�
|1�i���߯ �><��&���(���6��N�9'E<� ���_[y����~E�+�$]��vC^��h�]��S��c�Nm��b��⦊���.
�L쎔�i_p.�O�G!d}�VG����'O76
�r�ǆ�#.�֒��ZİfWOlq���Y�@v�0d{�y�O@,����h%Se��;����bM�l#���n[���ζ�!7�ۥ�P�u{mp��4,��lI���.�K�u%OB������J�!e��kM��z�]���+7����&Q��y����B�璂|������ﶬ@V��4̷1�ܰ�K��IU��b<��C���
�k���=6+�o�j��<B88����F���Unt�9��G��Z���ћD����/kd˸D�n�Ҕ���x`�,/v]�e�;�A�A ;�pV���������l�Q���V�Z����}���p6�̪��G�i(���?+XtI#���Q��`h�8܉r���yL���/m�����y�5)n������a�����UeQ�z���[L��m)����7BΦ�ˍõ�;��kp��!yZm3G�)���Z�^�g<3K?�%̓db����n9	�2��L���1a����c%Sd���J�4eƅ�n1�ȥ�1	'�0�~O���������r��=0n��� $-7�ſ�9����|R#Q�['�0�ʔ_[��!K�x��r�,P���]C��ɭF�[3[&�w�I�N��ii�*I�F&����<�y��'�3 CO�s�]5���3��ZIa}��69+�1bq�OB�5�'V��/��(B�yu���s��mO9��n~}ދ�����󙙊��3x;���_[��1����M1��:[k�H����̯�lU����>K�e�ˊ�F����A��<.�ض}�H^p�W��v�X�H�3+=	���f��k�tC�;Aɔ����V�g��E<��V�˒#�j�3Z֢��x�RةQ�k�Q��S���W�=m��\�j���~=W̓zf���p鬭'e���O�~�O{�73`�s�;>1��1�*g��/7��b��^��M�<yN	�/<�����祺�?�B�~h�g��Q%�����Ns�o�o�Q�(�~�!���/ːR�[:	'�=�`�(�r8Ӱ�:�(��I�͜]�C�QF�I�UM-Ua�M>���OJ]i���u*���I�Tp�d=	t�(Ő����G�$u �D��G���|���QX}�x�_�+��!��y����\!�0®(w�0�#.�-2qg��'�����%E�Li[3�>��t$� ��|~'ՄR����;�QlK^�u[:��5�ѭ�����P��GjZɓ�f�";}v�|�m�Pgt����)x�Cq;��w%�,��8��Gw%�q��8�zh�w����o��[u��1����e���ˁG�T�Ϧ6�G����"�]�y*M���y$��`l"wl��bϽ�t�J����L���d8�ia�!#3���=�'�?w��Mv����'z6=ƒɋ^�B%IH�8o�n�8)T��e
0)�E�C!`�^^UN(�?u#Ȍ5�
�_�rD	D���oJ����#���F�
�e_��4��3j峸������&��Djx�=#��p� pB�,��	f�_!����QXef.z3(C	��eD$�˴@֊ �,ZN��~�	6a�zh����������I>  ĕ������*40��Vi����?���f3�9�+KAG���ߣ>�Q}�6��~C}v<�J���U�����w,��������[�+J�H�/��o�Y[���kd_Y�/~��-�|���~dx=���U��W1c#n{�%
K$jE��9h�t<2Y'�WP��{�ﯡ����#A�)m��Eݲ-�-p��)a�X���f��|��	�/e�[�߁G�rt��Һ���E��y�{J��}~U[rw��hc��x�7~.����?��M�V��=��pM�����0e���l'T�<CH'h������u7F�<�W<�x��a��dҽ�㨫����*����T�IgED�J	J�AB��WE�.]:H�n�B�Dj� B%� ߹xyޟ�����br�̙s��:s��1}�4q�����C,1_.'���M<c�D2���Oπ��<�hae�)u����v ��IzL������F�4�)���_t��ȕD�}[�k�6�B!�T��&��/��;lQ�v�뗽�t�h�sS�ɯB�'���O\��7��&���������j�s6-A�Uo���u�7]Ώ�[a_�sq�:��d�8������Tu��W�&'��uՃ�Y�����m:�tr��w�:^�j���B��J}w$|���/O�c�����4t��� A���Fg�æGݻ��/���A�Y�B:���	?��Wsh�,���|�O����`���H���sv�ɨ$�$L����Zn�N�����H4�z�,WN�z �)�Yd��vEA؏gUg��ˍ-H��x7��tfp��$��_;qz�^�)��wS�[�rT��V�W	8"G�!��WF�w�(�@~�}�	�)����ʳ���Z ?O_�t�a'���e����*��1�c�-���.���r��}q2N|�}y~�(��Wq�Ni��Z����$#"�߼�0x�ks�i��F�0���^�T��]
*&\J�����he} �qif���K냫�d��f�.�.}�+�*k4ig�d*�l������ �VW�����M��k�E`7�l���h���S�	m'z~QTGN����]n�:���1r��@�@;���$�����_&ku�/���;�Π�ѽ���+�t�$oַ�����iD���c	�y��[�}x\	����瀃;+������K�����tWf?4��-�ҽ�YK��3�jc�x�s4�yo:��}�=�[W����E��l ��j`�:��W�a(:p���Rnя<��iW�*M6yi���MmE�;�n@�\� �H�q��\8K��S�C8l��U۷�Ǡ�z��ӉP��h�l���5��^�Y(r��F����Te]����K�0�Y?)m���^��率���9�i�ژ��뒮c�F������
^��sR�[iXOWX�Q0�b�/ϼ�p��G�l�?�Y\b������ �X����_�&��m�%H�����>+��}�jn�~V�~��F�3���(���D�C3��lu��$2խMER0AJ^+�ё�8o��U1t �`ݮa��:�穽�v�N�i�|e��閘���~�� �>�Ǌ���>�TK�T�����օ�t���s,Wi�.�ʯ�$�q0��o�����\W�n���1�?i�b����fg�Eq�!�����`��Ս�+\�::-δ�q���O��#k���v;�]t0�k�?������(l�0�O^����m��.�n���2864/�r�����TO�WM��Ik�w(���ۍ��[Zy�._���f��¡4�J��-��&�	��Y��������}��-a��{��,�T�`�ʶ�I?{��C�o�٫BNv_V���;A�}=l�%:w�`y3ñ��ŃJ��:���`g7���&���]gu����
v�>�+���F�j�<L�=�N�笛�lI��W�Rc�Е܃A�Zm��5B��v0��G��j� 8sY�x;t�%�������d��N@��.[���,0Q� �*�/�!��~���4��q��6úI��g�K��P�V���j/h���s=���^E�'���Z�GGc��gǬ)�/�F x|��_��馫�O��Ё�Og�o^�|�H�)+������2[1��D�i�;�0��J�*z���'���a,��	�{���0�m	c�[W���ͳ/𕚤�ؤ,-��cb8Ulg�Zk=}�%��,�N�n�����f	��Jo���\�ġ�@���0#�o}��/	^6��O
 r̚��V܂����#$�����ט�`�K�Jǎו^\��Y�rB��C�D��r�c��'���m�"�8�O�U�=��~ �#z���僸�o��@���8�;��d��&�^Ԋ�����=�᫝ʰ��G��v2k�[�9�� y����i�FBģf���(�����z}]��;r�X1阂ם�i�׀�!�*㈲���|�q�4"y�, l�����*����]LX�\~���m���N���_\����r@��p�}����`�HMǣ��M�J�*b�_��=F�+�%�Ux}��B��A �>JfGػ6ALJ�V��~��Ά�t��7TgGt͏�,�s�1)*]�\6��쫙 ̭���t��#�������A]Q4�8�W�Z[[u�k��ir��F�.�ww�$�;��a��e���l��w*�4�O��Rޕ���0-lQU��*?#�p����&��s�/5�^b��z�*3�K��w����
��T`�[��nV/ܧ�A� v�h��&��nv�U��Ȼ:�Up,`����k��
�Ba_]h=*�)���.~݀d��M�.�&|���Uu�\�����l���PX�����脌\���o��O�H��X\�Y���H<NCII	��y�^��5 8̚�����C�a7 ���u7�!���!7�zt���7�>�nf �y�+W#�3��rƭ�W/f's������'�åk�����uwC�p�~������)� 1���h�H�:�`�� �n�I"2�2~3������.#��I�����F�}�uٝ�q0�e����^<������g�3�4]��楤܄�v=~�a����d:L�c���$�R�%�;]G�p(!#�˥�pd31f�}�V��sY'�������L|X�j�z���ex��	�5-��&552}�m�tө@¼��6,�2q�M��b�~@�i�P�-;~�ڿx4�_F �M�������ć'��2,��f��=����O��[�׿�>x-CT7�������i2z�_8�z	�}%bB2Ew�7�y���/�B�����t@O���_�~7����/�k2�d=��=�dG�1�(@V6��T�f�B*an#��z9�/ߥ���K�v���l�G�\�"1��U�5*8.�3��r]��'��K:�W��Ƥ�>����S
�X4l�h�1�����1A;�g�\��<��7���߭ߍ����*�8��mᓓ���0y�\��*��ۛ�T+>(��(��Dy���,��o�%���/�U��]�p�x���L�G �x[������3"|�)"O�_�+�K{���8{�-�!)�"nk�����f*� h�f����@b��!mrL�srs�ʇ2���^��0�叽fݢ�4�)u��e���g"R�-f�~٫��/�X͔�|t��.�@��+j�#çt���l��wbw���l��]�56��2%��Zy��6��m+X�!�.8ő	 � ����T"3�U ����v�h���,D������3QQv���n`�{�v�Z�0�%�t���R���W9V.�V+x�Sz��h�nrҰhgsuvu2nX$�K[�c9,��左�Ʊ��u�ܟ�VR.�H���S���-f�'�.��-r!er�l��	���y��0��;��0���Μ��I�!7�̔�z�D�A77F�i
ރ�'��	�3��N���2�i�8�� �*Rw�������u���?���v��;�9�,��n<���3�#��}����M��������j5�����A9��=��C镕2j=&(����e�'O�퍔kv�P�[�w�JF�ok�yH^P*�땭�U˽��l�Y��V�TA���FJ�� �^���r�l��T��lݮnm�_Z�h��=��I=҄[F�� `��w}��t�J+@2#�~ -41�--
�X�U�T��=Y�Lqv6�ߧ�Ta��5B\�ș�����2���wGW�p�b����k6g�����]���q(B�Z@@@Tn��t�{ڠ�������]VTƴ^�7*��+6Rnkl/Hn����©]i�~Tn�=zר\���-�Q����+��Anm��!F:Z%��a��u�u]�y��jS��s���ع���>t7~��YZh�"��~�����ׂy�PƺI��(��|����S��Km^ړO-LML��X~!䀽�����cG^x�x~�I����b�6w}q��P�k��k��Ǐp�����|�W����p�P���A^ݼ�`����L�u�?�;������j�l_�җIN�oO�$|c����I4�8��SUHr�'��l�$��y��v�v��5�K+*��ߋ�PG��,�cW��_x��~�-�2¢�b([Օ�5�F�̸���W�a��sǋ�h����>hr,�U��=BO��oW`���S��<]���#��5�㘤��_��t�l =��,��}��GMb��^�_B�*(��j=�����jW`��l�;	]:t�s�V;&�J�Z@��}'�|E�T:������6��BH�|�h��H���s?cOz�i��1��N��!��R,? u�j@�w��uQ.�������yZ�Nۀٌ6�CF	����wc�nI�jvC�RK-�ε��w��Μ��9�̗�o���L5���|��<�4S��Wu�5�`e��
��VIl	������nܙ��cٴ����L�]��R F}�40�Rs���O�B~}1'ے*j���ZJ�=["W�Y����q�6n����v@u���s�����X ��ia�6�a��sNsC�}s��}������"l��=�	ٚ}���/�N�M�*���WӅ|��U�!��O^V��fp�&esR�������F�2����=,wLȯ���<�8mAI��H��B��V���w;0Dyg����D�ƣb����B�mo�pr&v�����q��
 zSb�A�5ͫ;<���z�5ވ�6�=x�?���[i����;v��Ы�S��(nA�o��: 7���I@�Mm��\����,����U���SG�Y)-�m[C��`��D���K�~0�4��^U�?���5����ra嚻�Q-�
�4��U*�����7��wxr䵝�+e���%1y�!�V\O����Q;��>v�baS}%ı,M`��c�ce��n|���o�K�fI��9+��|.�c��v�����M+G���d�Q���1����QMt���Px
���o��ǏM�q����	�����*/�R�J�M�x��@6�۰�%��Gq���3�'�YVM;5��LM��s��{.%�◫���m����7��ݎG;|��?����2v��������/ΛGZH>���K�3#ڪ��~lJjJ,��o�������M�p1�Ƿg��3��C�	N�Ya�jjj�%/�.��~l��b�7�����^iM����w������i�Q8=�� Μ0$^`��Z(��X��CIJH̛��ӓ�q���Č�dQ�)Uق������5�=��-i���KL T;�ʜR�;���>�V���1'i-?��9ױ���-�]�����f[48]�m��JI�KRF&a^k;@�«���3<%����Ro�����t�X\�{��i�A>1�O��>Й<�1�Lm�w{ǭ��-tAb\3ڄ�0��:�~��b�GI�j�d���+Ű��":���r$�&g�&���3����}_���c_�<������2�C^4Rhd��0Z�rH�YYΩW�d�6l�v�����k�}���V����[�W���݌d=wn*9lll�K����C�@7�,��PG �g����PKtu�ʞV�Yl!7MdD
(u"ѳ�I�M���YgX���H�L��I2������R����A�i����$�D�����O����=<u���rw��b��r�ތ�z�2b*	�	{	,p�|�WGKYU�����nŭ4�<Gk��j^�W��ѷ=,K�Okj�9�>!�7.Q�CZ��,&fI�)>5;�w��B&JT&g "�����8#m�ӥ90��߷z�����vR?�?��l�d��K̳H\2Z�j�튖p?��9�\�9�;#P�NK����D
b�(�v(t���O�GVo�^V1W\���l@Pv^�c*O�Y{H�����U��H��#+����&�v��?��{z"rz0�g�08_K�ʻ^ĳ�� u��z{���ߠ�$�
�Y[�Y��5T�*�}��5g:��1���{�т�ETy��m��X�$O,�آ%
*B������z��+�{=X�޸�5�@�#�]��9����1M֪��᠛}GϤf�_n���nOʳ|��Iq�-��Fջ��k��<�J�7q�
)�2_t^k�Q�u�L>��Qs7��c\N�0,;���궢�#!���#(I�p[o��Y()��Y����@�Ы.�x��{T�;�F�8��W��旡���H�J�b	�5�����V����沁)6�2W������Ħ]�e5R�K�����^�n	KHH zBtM|�%���פF��T�Y���E���%�B�0�����n�27b
�����D�!0I�h�O�[u,�ٻi��"��xc�ccxPni��t�Y:o���f��Uo��5�缵>��g?͡�\�8`�>Ojx1���>H�a6�[�e4��g�P3�0��JC�T&̆������n�qv���j[`�g�y6�|r�P�tn�v���c�o���F��mmm�-������<1�EV�D�q֑���D薾0�.6��w�	���9ۭ�`��;�nM���qF?=�g>��h�j�1�Y����yEb;��l�n�xתeE?�LtB�a�2�o�����<Gq)S��b�y�6�Ƹ�ZO�b�Ȩ_�ـ��SeQ�dM������kݏM��t�Y��L%Qk��M�?�8~B����x���M��}�._�������k=(��tmAtW�<������^�[��CԔm��ޞd�����p8�A~gɇ�Hj1���Xzmv���~9�<� ������*F�d�96�8&�ב�TΝ4J/�*/�7�>�E�V�U���m�Pߙ �U�TT��H��dG�F�m؂�h���짼��Uvf�^{[_��t��Z�7_-���O��������
�:����P�l%�J�����0�ø9]���dsP�p:p��� B[��sI�k��Q��ND�.����|\v�S<�p��� � �$3BC�aa�"O�dUеh��:Q�J��˞9�-��,�$B9��`c�a0z�;MU���j�jr�+��of��z/T�g���������'��j�8�2ǡX��������\��H��|%^v�)�����M��՟iF��f��C,���Ӥ�xd%W����D�(&9��_��qt��Y���#�n��R1��){v���g��g�%��<�;�ځ���%�[���LO�F�u����}�� ��I}L>�K��9�Y�0}&�>ǂ�p;��|��:;xHu[����e@9���{�,D0���
܈l*i��m��i�HGI���r8�6 �X�c���h%iQ�"U=q|&1z�ˑ*a�2�#��k#IP����*$Ȗ;+�K�pn�����X��$��T4��� W�����|@���H�=�"y 'ǥۅDs�>E�D��f�f� ��2����OU,d��* �	}4!9;^rh˾�v�0K��sń�2�)A����\�qn�:�dYru�n�����c����C�Y�'''�P1�<�����*Ae��^��:��^���IJ&	�M���w$\�&�%T�Z��^��K#V��oN�p��,�޾b��+�Br���5����1re���F.a�Rp��ׯ�'���}����.�c-�4ຘ�j�IbWӳjt[�J�0�;��T1Z�<���i�c�3���B#��%��g��6���b�61�D�]~Sk�����2T�c�<�������d��=��"4��Wi��R	؞X�<a�~�)l2�r�r���̝����»(�JR/���t�N&��3aD>t�`���}�*M�*L'���,4�"�y	~T�%Ҁ4��g��N���U��ER[[r��Ź�"��xi�F'H#ևܭ�k�}H���%�'�'�j}�L�G����.������Ġچ���\�o��b3x�X6z� Qߑ+if�~���sR���%:�[�+���M�g�JmZ��������3����h���pg��j�v~�r��'D�32�%���gڪ}��hI�����At�n�֤��eu�������f��sZ�:|Q�4�@��:{xH$3U�~�_�O&�15�����՜m���WϏ��;�����;��K��;�s�A����^�7��7����&T%
�j�7�6�%J�"e���l4�>W�\ (��a�!����nL?�U��/L%������e>��>Q&�{� �����j��lLgn\��E��*W�{6!�����Q]���\�P<;�F��ʫ���-����		�r�)�w�z������v޷���egr���928���Bvt�7�,l�����N��Α H�� 㪮����c(:�'�y�"L�xΐ��p��YU0�rdy>QhCE��c0��^t"���sۑ��)�tT�L�m�+qf�j�_f�G���v��_���u�z�D��I~H>�2����?Ҩ5`�N/����8�&����"g�;K��.!�kM�T�4Gls��u����B�l��T��lu5\���_��:m�d�"_S���>�qM�cKs�Q��۱�X|����J3��8�^Y����L��l$Q�`��؛?�R./;��������+r�y0~� �3�:Z�MK���e�>?|�p T�4��;U�WI���n��n'IH
U�����o���@ê�]NL?B�~�(Jd��s��_H�#�|=�B�%�v�Uk���?	'^Ř/�+����c�}�5���S��˟7dy�Xz�[���L<��1��GZ�>�%
�O����xK���/�;��2��{yRӲ�3��2�X�����x^nN"Ԭ3\�yˉ>��Xb�7%0��D��M��6���]i��V"z5T^znZ���^��k�I�┌�#�)�n��/p��m�>ݝ�6>$��iQ�~/�'��)�;��&�ؚ�qi���������Q��lZ��em���(�7����(��B=��zz윤����~	�r���n)����!m�1 �������$�wRs��R
��Z��J"W�&�g��� =���*KX񃒉�Dm�U�o�y�R�3����m5�zv����޳�4�4�U$}�=Z!��!T���N�$�7r��B,�Sv&J�J��́��ܩ~�uԽɉ��3���Lq9џ8|g0�9�3��9�_Bp��!��h�(�_��.�U�<� H�r#�̞0����Pl�Xt	�
��#� �Z(H������ezO۹@ �E�������/�=�F�w����d����=�3訛������,vR��i�~ߙ��CN1+J�oO �뻤]nX���@�n�q�AZ%PY����A�-:�v�{ڊ�x{�C�M!L��.i�
Kž6fä�
�o&�i�Ƨ��s�Y�`�p�\~�1�Y��iV�2��M�����!�"����hUM[��q���%�͇<�Q�.i�v��1]Q��!7*�����=�m���e��~Nq�����!cyL��*�e��p�DT���}�v�Dz�u4��Z�J��m�K�J�L>o/�	�V� ��1D[�t4��f�ϥ㻾ejm�+~��뗏B
�O��a�+J�<1[�i{��\d�揦����@�:�5܄ML������~@H�k� qpF�(
��i6t�w{7����C�M�1)��C�1�ZA�ҥ���i$Y	�e$����` ��3λ������F~v�E hb��B�8W&*8����ɛ|v�T��](99rR�n\zZf��*�2-������ĖIX]]��.x'9K5i0�i�2��DJ�D.m*��/Q0de���¯���`}��}v]X�Ў��'��Ǣ���͈�p��H�h�>]ZZ���Vjx��[�]�S��iI;q�hgυ"��O�~��_�
Z�z|��S��[�UhC���8OI9VD̸I�����_�]V*
D��Q �]<�p�����I����7P�o�#.Ck�@|� ����֖�9J�� �
.G���n��3��q��m�ȋ]�Qk�d�A5����~_�S;�h�_�'G�y�J�)���N�?��Bn&�K�}`�be)U�Bư�@�V&���[f�ʌ�p1��C�ǁ3%^s����PN�{��*�Xxi�j'��!�.��b7{��G��*ہf<�v4��`P����D��7���sϳǾf��v?��M�.K$:��5��,jbFn(J)�BR�J�&O<!ї۸�3t-�-dpQ� �ek!�`hf"j8=Չ�aQ׳�f��9����o�&�y��Y���&r7X���K6�ި�L6�;@���&	������eq �4��+�d(������=�j��9�u�%�r�}z쳆`K;���?�unv�k��t�s�kS�fu%jm	$�_�7��9��վ��JBpr[��.%�g@4�z���x���s��]���n�]������r���tc�12m��Y�M���74��툪7rq�A�慨@�)�mЂ@�k�� %
x%�����$�=l�R�-5��аˑ�Exࢷ'��^�	H1�5�rXڲhWwB�erҍX�a���nk���G�v[�(�"ۂ�fP��7��*�1R�~��1H��	�/��p�jB��� .�\o�z7��>&����GW�;��h���y�Ѿ��=Gk�����P/3s\����2 ��5�T�`'}����{�@��1~jƾ��0�*4?}��Q�u�\"d&X��;��{�C�N��,��a����4b��d��u���A�h �ZR��x�ڧ�<3LX0�L�`�{�D��� ��E~*M�G�4<�
ĵ) =6�T��ȹL]���z����v>��K���'�#��'�n���>��]ZU�K�Z�v��������ِ*�_�[1�t!�J� �W�r"�<�� �BYi�c
���� ��_Ly$�A�\���n�l���e�Ӫn���5Y0N�Ά�y��D;�Zk�C��`��p�Qe����	%e�0ݜ&�7��}>��վtJ_�mޜ5Zm�8�[s�����R�k��]����a��d�A���`�r[���W�\�P���k�K>6,.����h9KX������A���AG��lm��`��e%&�+�N�����M�_��k��= �	>���/��R�ݵkoM^;q�j�R�%� �A>�)��ùL}ِ�u`�Ì`zW�.�6LuxcP�O~�i��!����~gO�2�J_����_���}K=1�\FL�l��5q�p�bd�o����>;�n�~!��{�OM+����%@�^-Uh���OOl��VݏJm� � �)2�Fz��r�i��Z��@�2K��hW�#�I��׈(q&63�gg@��Ci8T�t�]_��"8ug l�"�W�	xD�f:Ż���3}����~���b鳪�$���8�f"�2N��	����g���þ�ЍA�P��]��i _- _���Y<��$ew�YŝWo���L���TG�ϖucD���d���1Q3�v�B��C��[�ò']��=K���2�r��0�ɐ��SjyL䄆(wWnGL��1u�� 1r�9�I%��3l�	{@)����A�ԎQ�/5��J�0��Y��#�!��p�Q���Hj���P��%i��#��v�y�v[��2dX�����1�S�%�T��7��ӏ�" [�nH���ڥ���^�pt,c�c�_,�`��Z�0�߳}y��`�;1w��������`K� �@�c��]9$J����7�`F���Wn�~m�"kl-���©�#hnY��#/�4�Ux�%��]S(���c -Or쬊��j��fE$��w�wŗY���A�&+>�,Rf�E�K�!���P�]�ҳ/xM�>'�F^�{�~�k��9uOɞ>�d]I4I؎o��x��9�V��ܮ�hS?|wd@�j�̶�k G}qB�8�Uj���L�q���#u�v�{\����C�˓�4P���ż����B�c����ӛ�x]h~.�`���J��2ွ��9$7�L�IL5��G��\�o���P��gj������z����l�c323�o�>����Jʒ\����˃��,��u��^�XN�W�K����?����h]S���x�Db(-K�ޡ�]<�=6�
�R�;52�ӚPB5�x��M�v�F�=�	�[I5(|��~o4��ȝ�Y�ԏ��.Yj��ww$��Y�?�>Z��Abqdgȑ+7o�z�r�ʩ�S�e�䆏Ys� �M�K&��ʇ唦Ծ�Lhn!ќ�y����~�5$	��a�Զ�x&//�e����ߗ�w�=e�K�f� ��S��1AMh�fPs`����f��~u�����,�>/ e`�U��5��S�3Fa\��wgg/���]���Dul�{~�X?�Ez�w�^����[E0�V����y8� �&X��DJ4�_1KF�ti==J� M{�յg�"�R^�V U���$lE��6�L
�>c~���H85=h1��[�'��*�v���t���n�z��)1 ) `R-��ٕ��^����Ԑ��Jנ��:hu}�_^�f1�BI91�m�x�0 CO���>U��^(��3lԽ��=����{ȄNCeee��l-�Ђ�;�b6X��J�O;[O��h�ĭ�<X^.S�'����&���E6p��ԑ.#�3&�s	��Op�g>-���~��a�("�;���9��Ώ/M��i{{o�����a;��ڑ�F��_���x�N�Ўd�e��U:��8�E�)��8������%����9���>D��L�є�&'>�ݰ�8�M�X���?��)���>��*.f���E�j�!�BU�۟��B�s1yh8��ں� ��i�y�~SR~z���lR�`���ZLڝ�/�����#- ���1���c�N�-�&nL��dк����\�>R5�g9<����Nd�]�:���	R���rMu�H�4,�s������q2^��#I�i�~�}�gM0�#������+��+����$ƍ���줌���$���$l$���i!@���#�� = 6��Q:r������^I��l�{��r�G���J�Ԥ5����[|�q���m�2���	���B�a�%�ZX(Q��٦�ZPe)��E�!��r3_�i9%U�Zj6�/)od3���`pw���X�^pl�	��]��Y�5#�6�E����S<w��w��I[��[�V���S72
�����ho�=�� ϗ3�:�>�\s��b󦰔T~�_Ϡ5$�"8�+�X�~���|�E�?����������~2^���3z��N�6�Ա��O��u��)����}Z�P�>��la�p��Z�m�_�֟b�e�h���i/���+���=�ӥ �ձb:#�,���j�{zM�<�������}��x.����������N�6����rˡ�Ko᭵�
�OlS���NF�Ğ�[���g'����w�����[VWW����T�P�ؼ�|���2C��93��b����j�)��//���_�K:_NMM�qtDC���\��_<����<�Vbr��X���1��y9�/9E�-.:%�u6���Pմ%b���ǖ�W�dWu���9M����*o1�U��x��2�fFʩ���5F�Ц�A��e�8!�;RiʯE��{�D� p>���Ǐ�~�r�$R���	�i��`���xt���ϗ1&o�~-t��z��I4�}6D~ǃ�¿��!�Q�2��3gơf�"�n_������x��:��%�� ͈s�j�&���Y�?/�'Y�S�b(���+p�o��bdG��J���]��,r�(>"��W�[|<Ж$��Bq�c�'�r��o�����6R�<)�V���DT����P�[z�`1�$~2���	,ԸE�W8MX��ʊ�@ٮ�<;D,��]#�`�������vh�yx��ٹ�i�{����}�:ٜ��!�C�6�
.��������x�w���#��j���!�nZ_��YS�{}_��Q0Ǧ�r��sz5�ݤr���u�}mv5�5,'�Wrsrr���������oZ&�d������]?ʺ�|���+!�T,���:��{i�s��暍:�=X�`)�Ơq����|�N%5Q��=[�3��[��1L� �);�V���_�
VI��[Db�-o��5hK�nN�ᄁ�������J�?��.l�&_�c���V�c|���^n��W+��S��|z�S�����O�Є?c�����7qD������y��ښ�c��K������A쟘c�Ρ	8e�lu�W'�*���P��B��FȢI���#��g�D���sFf ���l�v|�9O��6���W�!�����Ib���9&۶����-͏ݶ;��K|yy9vn��3�rC��{526>�׿�"F�RCz&����D�{�*�;y2�u���$˓�/���IzW���P6i��9�}WR$+�{�YZ	W�XZa��M��ua�w��ӱ�/~-t��kmU_#�~�ɨ��D��������:a?2�f���\�k��wM�ϐ�l�;%���6!���4T$XLRo_aE<�G�"ot�/_�E�Z�aº A9������2Qr?�������L����+�w�ݨ��_l��L��ƯV�Eb��}=8�x�=\����Ɩ�����? R��{��PNX|n��z_�	ԶV�t���3���}C�b8t�ѭ'�Sy��4�CD�o?��#���-�Ժ*�u��ω������=�^yJfF�X/g��s����3������@9\~Z'�����l�s�(;���g�r����n`u��]�=Z��gBR�v��">��;�ŋTA���l��9!v�0���������7����:㊀��+�@�J,C���o��e�c@Q#��������
���CX�tss{�Ƹ/t�@7��L��4�Ғ	moo
���6���
1����Dg��eA�_A�����M2��Aj�������j��&��}���`����6�&���)t�ٙ��N]�W��_u�x�S���N��ǹ�Mb��_���=5�.�����'롽� ��ȉ0(�����q���=�mT��l��`f�J�����������7�7��M-Sk)�a��O��&���L��(ݳc�I�܂G�����t��7(}�΍�3E�Q��V'�C��Vg��?�x�����߳�`>m`�������|�՝xƄ;��w����.�*��/}s:1�&�J[��C'���U&�-�|j����$���-4��.�&1j��$T��"~�Z���� h���ׯ��d��A�0��������à��\g��.`��J����x��s�j�c��v4swr���ޛ�:t���5�#Ф=������ç/�@�����m;-����ĝ���k��'55�������-����5�;_g�?�K����x�l��E�MGG��򣽯�
=A�D�|kLY�UR+���+���P|�W��v����m���,�@����s/r����KK�ߌ'�BB^���W��-$��Y��K�|���:��g��mq�/����;a�J�c0��7U 7bqm>i�z��V��m���Ǯw����Y����A%ї�0~��k��7W�L�X�����O��9wmVY~�tO�^jﶣ ����/���DT��� ��D��Ɍ��#��D��Ћ��u�Y:34Zl�A�r���M�IЇ5u�;ߡ\����C�l�������Dog���_/#PәI��,O�\�u'$�Ͳצ����\�4\b|��'3�.l�m����w8�]pCT	N��:��KKK�L�G�~��&bkg�&�3�*٦`��O���,|_e�5'g5W�E�z�U��v�%�x]��}P�K�_��.���@��zz&Eµ������dÉ���6��Z�^r��%op�6R(��|lx�LF�0��� ~�DO˹j2A��}_T�!�6S�1~@�/E21��zK.h�G���Q�|�c��@M �m�Y%�}��db��������3)�?�31�0!5�]�l�����?��ά�HWCD=�����x�����w��U��Id#]]�	~E�xori"\k��P_�+���`6ր� Iכֿ%I�,`f%++�|� /��{��	�,�)��\^^^�>CF����Yl�`�>��u5G�Y٪i���T��Y���+l`���'h6@����9���]���R��Ĺg����M��K_�C��?;=�Z�l��SK^{-��zŷ��Z8�bVʌ�~-�E�K�@\k����V##�y6������eα��Xz�$i�����h�]J9|�k5Z���=�}N�}��J���b�I���O�س�9�s�عf��3U����;5�kB'�6F���G|��A�6����-%&���A�8Yq��3�m�����X�ǻ{J�(��o1>�"�q����*�	��F�0�	d�����=~ iA�������n��l^QH{�T_6�����m����� �:߀l
����=ON^��4�<8������g��&�HRϙ�!��0�#/D��zoL}x���0�����`�����o�>�z��{�	�@g�]`�A5V`@����|f iu=�l
�R�
w]�������fw�@q^K��;e����ډʴ禪�N�8*�!�c8r��`�%��o,Z�pR������YqQ�Q���8�[�%��Z�3X�w�����2�����|m��%j���	m"S���o�� ��O��h)>&ÈY������к��f�/�:��F>�8
2����ӯ���,~1R��r�[�i�z�ީ�����RGs
�?�>�砼-��mA��:�/���Lp3�7��1��Cj1	�^���k� e�:66�����:�
�s�#~��`8��ܬ	�ZzA��������ռ��#~��Ǎ����	�>�9[ gyo��|�]�OS	wf{vq��օILR�,��ٽ*�z�T0^����>�c�~F�(|��އ(��	cu��\B����g ��r��l�^�v�)�\���б:#�-�դɍ~lux��<�&ծ��2+?��
LPI������o����+-{/�]���3p�Ԑ�Sb6>RFd��D�]Me��/Іn�����b{__�,��zVxP��j��c�ɞt<2�J�����u1V��r7�mbO���y�;�{�u(�j�w� Ғ�A���!P�	:?�E�F{���?����9(v������,o��Ю��dA�S1���o������rR�&Ɂo|4���c��Ӽ��Ҩ6vV+�k�H���
Y�.���"s��8	���@�[�B�g�
���{ �C��x�,�F�݋g��wQ=_����ZK)��D.���Q��� �@���)/��:h�@x��]ڮ��Af��-�^��؋�m��4��c�f>����.���l�!_���c�����F�������
L����l���W'u�2#���3^����Ϸ��_�5<�X�m���5v��w�3���".�Q�͡�I#����Ng��`/Pv�p&�����+�a�Q�sy/}N�i��������1R~��S�6���J~/r�VF�3Pô9
l�/K��8���j�b/R*��Z����BK���S�lu�v����]T7�2(-�{�0��J��g�9�ˑ.�A�������H��Zp��J�p)l��GL@�e�>��P�{���u4�8��B�ޛKX<l�'�u�������{�yAMT�ݺz��M���۳)E��#;�Y�x�u�z;���x���T�O3�zG���o���z2WP^��C�	��=�q���>�։��ڒ%�'��t��68 �u��e��rj��ݾה�
�Tʣ�6@���w����dojY������"�+����D����|�.u˫	K!�l�=�8�=�*9�����dT�9���Ç���l��AOG��m�W���i4�)i��S�W"�T�]M���������۬y�V��.��(�S]"��[(��8��޻���B��2��$I��BZ�Z+���JTō�����fi�T��I8��H���?I���P��Ɠ���c�-��Z��a�(�@DB�CZi�nPRZrhT��n�$��A%F�`e�a�n��������%�x�l�X�^������31BJ$���ƽ��Hg��������I[�7%�掸�`�_8��Ғ�#�� �r��4�	�b;�~x8(7)����Z��V�O��:�_s��!11W�>�Uu��l�c��t��;��*ãS<�Ӛ���5�'4��^�ϾS���'�f}��R
ibg��s���	vR�����L� 	�[!;��J��I
�Vήf��I�S_�ǝ�D�vUf���	��h�����j��u������h��6h���e���D��r�F[�C���5nv����J�%���)�p�(�2�8"��/M[?>�"Sd*q?_b{�,T�ض������ez�(H�>?��Y6��]�����r���O8?�� ���Kxjr�bǓ'߂�an�U����,����gv�4���q�~[R��R��q�����9wt n�܏�q����Z�6�֒��y�>�~ڸ����R�;+�{ �F�x�P�J�>2ho:[�2���f��ô�:��2c�E�F*	83�l{3��M���ن1&�u�7�WQ��E	Ѻ19� �v�׈F��%���'�[D��sz�ģN' |�ǛZt8:c��c�v���`�N?�;ڽvҢj�S����E�=���g= u�Je�8�Ѡ�&�Q�-�E��&�ə�o�{��;��QY�����������W��X��=׈#�X�L#F��L���0E:��������.���M�4���']ϩ��.or0<������(�!�c�-�m?���C�nh�{�6p	�y�?��Ъt��g������4�ӇL��O���ޙm����^,��zt�joNu[U�a1$��{+�uz�	)5�N{��(����M�<�ڐ���{�ȇLy� q��z��׿����UD�X�{L�"��JA��v%7�G��]��gk*�DM�Q��="%d
~���s��9�ۘ�e�п�����f`���O =$%##S��61�v�}�Ȇ�� � ����KQ�eq1bfo���v�}�~��4?[GvEF�~��`~n2B�9���`�8Uؓ�7�uDb��z�i ��	�KU_7-����\U����Y�|�y ڋdfa�ilBrqW9-t�6����qm]ݢХYc�L�}ι8R��@�`����a������|> 	*}�t����;.Bs;���c`t�ifؼq)�fv���(
���}bbuky�L,��)u��b�Pr9�Z��[��rN��iWTD^�A&ehhX�cf�4���̼�3���6�Z;vȸ<�N��Z���w���j���yh����V�O��P�r��)�)λ�)ej�^��Y{��$��S�z٭4�J�O���Ylqvm�m��� % 1Z�>���aIU!���U��8�L&����->�f�(�����ZV~�z���hl�]����n%��V�<p]Hl��W��o4xeh��P��{Tફn"���P�� ��g�g�j�K��-���3:�Z'P���[:�6y���T�2���[�D"����Y��e��T�yWtu1>��TB�H�Z3��x�"O��� Gy�:aZR�?8�
�ѫ��7��y ��Y!&��������>GGJ��陑E��	c�6��}	Q��C{��=ʢ A�@QeUK��t���9^�2A%O:����`��FL����/�	Z�h�͝�یfES'���rt ��G9��Xc��) .&�ieo_ ����n�b�'��9�~����sw8,~����O����@N�tG����x���Լ��\�cߓ��i����r�����e�|�h���5�&����?�F���<�Ydu�-bS�ڬR�yU�E�η�!��PY��^F���}s�~1�op:U���f-�c��Q�!�qYa/����(eb��_u0O��L_D}1��T2�ݑV@�-�MDI<�0d~���M�"?�Y
@��X�eȠb��C��a�H���I��;�>�bAL��d	_U�����k^�4h��ǁ��n���f~$��{�I��7լ8�ޚ�z�:����P�~E�=���[J�~�vb6P��dԘ���Ϙ̵�r:7���}`�흾F�(�_��8A�cp�QU�����[������U��-�j���!��0��m��$��<q�`���Y }��cP��sw���:y����1�i��nM60�'�+pA���@X��e5&^���[���(B��ZG�yQ��'�x�rRטXe������i�ǯ�r����ȁ�4w�g=��p=j��a8JC~d�kk�b���"���&��pj�%�r����;��1?֓��z�t�A�ᾊ�L]o:L&����K�1��22���"K�x$���� ��Xf����d�	����>.�|���39K�%>+W�&�����sG�9��]����b(Z��C�]�F��(R�C/�U_�W�wˤ�I�3}n�l��t~f���S��\[pCĥ�g���{2��:���Q�Q]2I"/gba����Δо���P}�qC2j���I�HE�e���_�ϳ'7Ż��͠��T�b@3jz�'_"��୮ep;3U@� ��;��o�+�l�]�sI2E�o��1-:�-Y�F�<����x��z�w���Y�����+�_-���0�$�2H�����SE���mk[\��k�Gշf�9�yл5u���' f����b�k�u��^ . �1�ǭ�t��}�Խ1��A���b����Z������x��aYCS��ȟ��IV�/�ml���K����+{��~�]���ѕ���%!�y>4~�T}�\���kZD�,�d������I UX��*a^�q8��}d$)����8e|�c�VYBO�g� �v�|'��t��s H\^�ZT0�G�FJ���gK��l���:��'�I�q��>����95���Z�4>�Lm��(U>�q��X����~8�rq�ā�q�ԉq��jE��bӠ�¿�}�Şd.����x�v��r�������DR����N_eϜ�b�������j/VVM_�X�X~�������8#�F�1}�楩��M�	��B�Yu�ɯ��@�ڢ�r�����s��6Ͷ_&��AV�Vվ�O�ݴ�k`�٤���)��X��A+��0z�Q�0P��^H1H.;�Ś�"����p�oT������2�,�%���3�p�			uI^�|sx����ŕ݌X��7��'��F��� *q��e/ʟu��$�)))�VK*h���Q�?��P���=|E �kf���[GK����&�oR��î�9⹶�|m7*�a; �J�9��n�z��"�3�/c!5�0-�j�c�®1���U�'{�P_|(5{��x�����r|�Q�[��H}R�A�jj���У�Y؋ч�ɴ�����J_E����+�Ȫ{�v�+@9���2@����^\��e�7_U�u�S�f��Alg�����G]Ǥ�4E�������3�{o��M����-���/%E�wVd5jGzƚ�9��~8,f n�*Z�/�`@�<ذ����	��N~{z��(z�}�<��$�z��>��%u���G���D�ywBi��#˳h�ޑ7�*�ɢ���T�%1�4�ш�׷_W�1�E�lQji#F����?M�R�S�ǡsr~<80p[��Usdl��5��	�7o΁�=V����U�®��8@
|���pK�%&�;�cR��j���w��ܷpʪWG��9�/�R�I�]�w��\4) `ғ).��:LTуY;�F���ր��Y�r%�N	7ܑ��D����<٥�P�i�J����R�Nzw��.�1�ҍ��ߜ�=�j���0�����Ӎ��z��7ڞU!��3Ծ�%�4��I���V1��N�SSt�bdL�F�s�װ�
�7@V�l`4���H77p|~���inV��r��jaYY�P�vE:R\p�����7�2�_�jip�U9�@�Q�� ���yʗs��=<1MN�#���e���<���_W}�ǘ��z���K��&�^"��
��;�Bd����JL��$
9M���὆g��p�n����l �)���t�� u����~�#���Y�E��'�%�PMs�S�u���$"b��tB��::�Vۘ��y��Wu��*sU�;��_Q�ٳU8�S���_�3?�:�LQ�w���f��[-�e����p�ˢ?�zs�?�	��kz<�vXR �jW��X����Z�=,--]�,v9�Ϫ������FZi��S�kԕ������i��8x�*�FOhb;o-�荎���f��	��n�7�X�Fu��,])J�)V��i:��{ї1��|�}:��f��$ <a:�͌n��h�Ff�"����~�L����d�+���`���@���T7��|H=7��ֹ��@����`���v��~&��{���Ily�7hSGً�b?K�u*7�js��b��ʷ��LMm�?�WP�'�����`���\�H�Rǟ�|x���69�J�a�E���u:��1��Rq�g}f��xy�F��ӷ������<W�����JJJ P8o#[�D���W:�=]j[H4���˫��
$��������:ӏ����s#�1P��!���/�6��y�X��D��u=��_���IUu�Zf��?�����F��z��X$2ڼ��쨸%b@^��V����*ւ3x���nP��Ou:�
���[�RǨjh��yN��@��Z���߳,��X���c;���*�?�:Ψ������*�������3F$sq���F&�@t�kfM(�*�s_�m0�ݏ�`���s��jȔ^���R�JEm?[����8���7��j�"��6,��!"�6ߊ�.�Gg���_�ڂ������kX� ii�$w�b������"OfpWW���&�}S��Q����,�������H����R9�r!�t�,Q�bH�!:�����K�M��4Īz�e����7������\G;��ҪY�B/�#p����jq!*-�z����΋H8�z3D��Xu���Q�+.޿n��X��
�°v��2hG���2��:6GT�$��n�����	�?;��r?F�1s�>� �Pr��9���V��'n*� �*����B��į�Ƴ~v��I��N��d��}�� ����G�m�L�x�* O����yI��⃃�$q?�1�}dP��F7,�=2��M5��BHKKwTG�,'�X*_*�qŸ��1��ҟ3/�S^޹�BJ���փb�'Rֲ[q�ס�Ii"���IjY�������@��2)g����mR��i���V�3�)F���ƿŢ?����,�8]�V��}����_D��[��n(����
W�\Q56������]�Z���� �*�F��&Ʉ�Hj�A�՚͞�p��>�ȵ�-|�U���>�R����NV�x��MC��ڳ0-~B\��Q3�5�a�3����-���O4��������^�"��g�* 8��{o��:P9������9�'��P0�>��n���7��8�I�[���5���W%vd� ��Y*�]�d�p�ٗ�R$�;=lr�1�c�3��d�&�	St!�@�/J[�#8���N�#��aSX���R�1�4"%$����OM^~��%���(Ak��H�R�=s�,�B��'���U��
RT�}y@�)h+�3�%�G���ְ�Cw�R��H���uy��؟���+�%��F^�y�;���:82ZVB�����{�}�M�q�}����{X��ֽ%�����ǋ�~��C^Z�݃��j<��	L��$��D:eV�}ܶ�5�E J"�I�A�w�GG�	����|��̌ ��:���)R�ݳ*jB`��G��!�<�Yt[2���S�i���`'/x���Ȳ�����Y�6#�FD\H�O�DO��r	=��Ron�J(:���l/^�fXXs?��%�mK��>-�P=aa
��)
/�g\��=��猈��X����)�̥�T_3��{{;�j�C+�-�QD�����*bɘ{W��� ʦ��V,�:�{1ϛ:��`s<!T0�N��{���A���¢W�����2̤g�E�$&���� �;���F���nX�F�'�7�8���y+�{`o��?0��Ŧ7�����uMG|�/2�NǾ/!y������F��Gg�, `4��(e�Ȯ���~g��͛;�U����6��<Ɵl:���T֑���S��H�x�9n�iX��JB�ɵ�E#R����}[! �v�--�ka�,�AJ\@��4$�C�����F����`QN��M���{���}11I��XQ5�Ð�^i W@�����:�����	��?�ݺn�a���rcnsӢ;:v��4����� #u:|�Y�H��I:Ea�7�5�K�|9��?(�2���,1J�J�#sy��,�@;i���g����6a7��<)N��bc��m��|A1׽�=��%0��,����qS�
;f4��:(����Q��=7b�M��M�s��ْ�J�r�g�6�y�=��R�6W}�ً_�זҎ��j�g�rr��{��AY�n#�N��wfj+�xn�1w]G�*�])�%O2饙�Z'�#��RO�_K,�?Ο����Z0yJ�3`�`6a����R���8&S� �T	�1��מ$�؉+	g!"���Az;�{[:��
׊ .�.�djsK�b�O��I<�6w�e�1&-q1�|.������"��E>G�g'�5�^��]�����q.M�mA� 
ԕ�'�O����s���>�2|����0pq���^&��(�����9��T�Qq_�V���ͳZ^�W���(�]����lu_{���T9���mC:��� LP�F>��ԸH��W����RP�i�RJ�^�tD�����o`7��0�Ŷ�`���i+�\٦�Ŗ����DT�"J�#��g�v
��~
FЬ��SO�7���i:z�'�����σn �-Q�L�/�UX�b�M>I�)F�m׎L�@)���N��{��(m�=�7��0������ �����{[���^�!����8����1�u���Z�!�J��׵�w�&�.bfo�:��ڂ����jĕH�x�td_�
�����\C}i`�D�Z
˘#n,��w�|+PE�"W��N�R�>a�o�:c ys�J��	����M��/A/ ���6�p�0JZ�>��H?	a,���hGy��N�c9B����W����>��QSˎ�ᘖ'�k�r�"��b ��Ɍf�E�޷`g�O�*�>z�LN؛RIhOY�f8޼=_%��V�����gw�<l1IÇA���#�=4l T�K�3)x̲�N��x���[�;�� 4w�v��Pg�$���:S��8�֍�ⲴB,�)�_K�Ư ]W��>/߭���aT�l��h{�9��]�|s�5��Զ�������Q�D��a2�}2�{#�8��a���Jwf��t�Xa̵c��X]Yi0x����M􈾰"���L�~��!X=��H���>ث��8���NO׎�iG��ζ�s��lz�~t��hO�q�x�dro�/#��c�|��v,vҋ�t�"�)��~�ˡ�co�~;@3M�"�2�pp]��wg�Z~]�[fs�m@�%S��Α�^� ;�p��ώ�7������H4]����O�*��OL���GKs�zp�PΦ��r_�����ѿ�H���h9����t;�ݏ�5�֚5��?N��Z,,�;�Y����`�A��`Tb��s���P(rr�H^ӹ��'��G���Ҍ����������!��	����|��}��[�Ǽ�ϭ���yr��/��S�g�hٙ���G��,D����x97D�r���9�h�R@����ʶ���D���d*�A���P�	�Ԫ�Ō;�J��NX��Jk��.h��Ѹ��G�4^�[SEWhK�ۨ�E�����Z��C���	jg��% ��46[�����="�(%M";�,��t�{��6�%��ԛ�
�Z�����SIS�� ;1u~n��L������|���v|�qYHmjL����c�yۥ�85�X���Ό�ω_��ƕ]�K����E��b�9B@��It�`�!J�3+�Z�٪���:��vr{=2�[_�}�gjUE&v��7=���`ԯ��Sw���m����5:��2�syQ`�@	.��چ�	�5b�S���|,.���dRn8�t����7T2�"�}lKM"�j�wR8h�ݜ�v��w�f|7������
�v�M� q�!C�ȦT�;G$�͞,�V6�g�xVV�B�����i��k�͡����- �p��=B�Q��mG�>�S�F���8-t=������q������Fjq�B&����=|�X{B��B;��C�(�v��L���]����Px�������R�/�:Bh��N���4��	B���|0`�<���-��p0����C��T���gU�_Y�8�T�[�GM��	� �q�5��R��e3�f�p�r0��K4�Mҝi��B�p(N#�6+���?:3J.���'�m�&x�`p"�`VW%�,n&oຑ&h��2��_v� ���sOXv~a�G�����P:26��[�c��>_��aQ�]��_2��T�`�iS �O�x�����ҥ�Xuf��[�뙢u�k�@@þ�����χ=��)S�Į��N��>z�ZQP$-7}���Hu�hB)v���_]C� �Hi.7��/T.�����7
*��{cWυ;w0�'����<��+�R�Z����+�=�7����Q"|'� )�Y��O�(�2М��3}����-ο{��N]'�=C���)�.H$m}��5U��k�N��G붎�W#:>Ɍ��~_��͸xo/�ģd� k�bu�F��&T��Os�2Q ��r���`тO���������
�6_�2K�bK�=nu�2���S�)�̣�P�N;���q��Tf��f��Ju57=�=�Z*  ���% �:8Hae<;�gt�&�������Ӯ�m��-2�����K�꣭"�Ƅ\�~�=)��N����+
��kt��� g�������_��֥�рI��H����V��t�c[���XQ��{>�r��so���"N{���A�~��`sZ�Gc���9+'��Wq{�p˵��⪤�l٫�?u����Rlp���R-�WC��.���gD�BnĲA!.��8"�ԶP��紜�c�
��k:L=�m2p
v#!�~�Gb�@0pਣ��9m)X����Խ��}Z�'7~eC�XD��N`�f�J�R�bRե�����d[�=�cj�<��sJ-Z p0m���[U��:��>5��Fn(~���s����(b�/�7�Yv�����ʆN�7}dŀ ��'��&��t1���́{��7�O`���ut��ć�ڤ�⯕���$��$��e�[�6Q�C 7v��h#�YR����C�X���J�^��[)'~��`q�閦�����$��qI�� �x��O6�l��ޞ��&����������$$P׭�rT�A���������£tܘ�OTٰ�h]�SQX�h_�k+�ŅJw%g��S��LAFe��j�L��r���;2+��_��������S[?�e�Jkz���z'� hd������?Ƅ	��6Oe�i�uVy����p�KPVZ:������5IB�(5�ٹ��X�]�Q,��O��82YC-�k�R�&�dɲ>�N2X�{��/eq�I��&��b�ٙ�ڮ����d��p/��)��1��Ȏ5���]j���������'pW�#�~�)m'��]s��QLg2$��E[D�Ţc�. ��'4�<CП~�d��� �$0e����%�P���.���������Z�4U�� v�l�P��y��
�H��zr����F���\��HM��������7����F@L^G𗋙���B�q��f���x]��1ѷ�������|*"%�	]�6�	�K�"�G�:n�$.m0F$�ߕ�4�r��'��a�����<ap	��M���B�>����!���n����g��om���6�o��c�=�u��ZХ���vR��m}��:���J�6��z{gG��
/r��IК�C��;�܇G'_��H]z:֑��}�"it�fi���w�)�=c7(K��>���E%�jLU�)j''��Lw:ĭ��`06f��A/����N����V�)���)+�-�$7LoK��>�~a�BWs�=zR����✱i�
Qy����[�u�u�j�U�+��ؘ����j�|?�T�p�}_"��~}���yqY�O5;썍G�_ŷ�Z�y��˥C�"���Љ\���&L�jXeǼ��� Z�e��O%��ً�)���4]M܄ogz��2��*��B^F�Q�GU���f&>y.;�F*nM=��8*j���\b��ܸ�`}�[%��M�K��*�����1m�0m��O��ѓ���;�:A����g9�����d:��G�� r�`�����]�[�4��U�������ħ.=>%*�R|lF�c2k�I1e(�`�Øۡ,O����W7��Kc+��BK�@6|�����c���d���o�Ag����^ǹ�y_=Q�Α�m�)��eC�=��rx��V@��'Y�����=GW���,]�/�Ƙ)�����t]�`;��<_��|��_G�h��B[=�/��8�y�h��ܢ��W�uq��<�R�*�}���c�$+�g�͸V�0�@�N�shDau\�6�8�
�?#fD���0ߋ�6�Rs��H�D΅*�T��G¼4��s���rBZ���ߍ)N�Q�ׇ�ifq�35Z(g(S�K�LT:p�P<��wh���ܨ������҅��,��{�s�������:�|b��YxOJG�l^���Pl'#�}�(�t�J_!n6�-��Қ]�0���Ⱥ`y�x��v�^����ʗm+�.�1b�2����������Q��K��ڋ?�j![?R���ew�/���s�q�,�e��-hZs�s~�*�t-��1�Â���O=�T{�|���7ښ���sA�7U�G�7y9�����:��}�}��8�f��3<j��ZE5���~-N��w�����&��$#s,[�,W�d��9!�/�7݊��&E�a��JM�Mff��V�q��R�X���骩Ň� ��\1O�Ǆ[nI�g��y�L�[��X�Y!��+����Ww�����tT��������u��s�Q��x��u�T��A4H�3�Y�(��=��o%l����_����<%�.nC����w��h"�B����t��۫�dl��\e�f��d�����ܙ�����sZ�=0����[�����|o2>T0�M��;��&�����M��F�<���[�,�7�K��Vo�U�2�|�]����l-֛��BP{�����ׅ��9y����uܺ���6wfz�)n�efw�Ruzmơ�i�Vj�t�` R�jd�~�:a��D>���O	�ͮ�3���Z�c�o�������ش�%ZD�!�y65�(ҙf;�,��r�����J��Ρ"k_^�k���F���u��빋~��s}�M�"q��r��	���M��-ɏTފ��Kb�\��IU!�������O�G�z_�����J�Z�V�!S��	`r8�r�t���&��>���Q�ⵆ1;H7�@��*�w��S?Ǩ�����I"{:����Uu�f1}�R�tM�j=�S3�Fh����yi�RC���K�};Aoܺ<|!����
��N���p)#%�ӰS|�IpפU'�z�;]�I���f�XEo���f���W��!N����$���m�;2q�,�!|o\z_0��k�>��c�tLR�����̠�U���E�xawi`~S����T�Db��X�]�Ӽ	Y��v��L�:wX���mw-���dɱCNQ�� 4�(��h�.�ޠL�W���O���z�+R�u����ǖN.!��"-����"l2�e�5����B��E����ۼ�k��-�G��+ۡ��9�:2+�3Sc��j�*�)�ft?ģq�|Ol�[2�on��߂���x�@�K4<��1��=z�l2~''��
����@�J����cv�o*^��7~��ϻ�8K=RE��z�+(�XN\�@�ȷD�^�]��E�O$�8χ��I���;@D���y�����4������u�e�8�8�xꕯ�u5��\����Z�1��q���\�-��Y`�-eZ2(U}����]$��~lU��ܑ���7�wN�F;�9�p�7L]���<=�l��3�J�8Y��Y%�)_@�v�'Ox�?x�b��{����c����P�t$��]���ꜚ��T\?kI��]�zv�m�E�<��T�P8�dd&�^r�` �χ���2M���6Ui���[�n���R6�e�ܓ�e�Þ�A��'�L	M���$h��m��l�D�_��;Z�q���\ȳ�͍g���A3ߏ|6��A��Oğ3_�;�n��IcT��a�k�:�C�a?���YxkY�����.����Է��*/����P,��p�w�n���TBq*�~�ˤ7��c���C�Zf)�)r�����g����i���{!��a{�Ÿl���E�v͕)��~8����Q6��7��>��j��IO�}�(��u��|�Q��wo�Qu �(��xu��lvi���2���������q/BϕV�O�#�� R-S3C+H�~�U	�X���3QT#��Z�P���������>�"؞h��V����n �R���$�[�����:�����92���yC"M��%�9C9U�rC ��ڹ��a�9�4�lyk� N�qB6W�	�'�E�x޹zMn���P�B�*+�k�ە�P$�(�i���2�>5iN��ԟ�"�t�9U���u�"��r v\�G�(���[cv��w,R\!N'�z]{� #ڸ�n}�V�Q�33��f�����S�.elќo2>`�e�����ə����RTh��Y#3���
 g@���D�l
�55���s�"j��(�t�՟��4�ҵ�����V���e��MIyZ|�SSn��>	H8��2�� �z��sv5^`+����E�}S.]��N8{��Tǖۃ17m&�1��Ѐ��������}����+i�d!t���A�[���?v����[���,�x>�w�x�OOƪ��|t���b@yRrI6�~�c��n�M��- W=��� �ql\y>�T(�X���R��zZUV|zAY֮D{�E-g�*� g%
2_9|�"MB1`�'87ѓ��:���:bn5�Ftճ.%���f���Dd(�m1��^a^S�F���?�a6���i���z���X7-_wo?�2Ά���<@���]����y������W�b@���s��K�+�@U`[�c�D��,P��z��&%L-o�>6Z�8}����Yf�����7|�|`K���Y ��o�1���Qr�9�/b�2<�۲?��_��rQTn��d�o��3��`���ӌ�ƲJdQ �n�(y�؄�?9���V�y8��RiCz>�#�3�����?����%Z�#���8��3*��i
xm�zz�P��� �z�I�j���Wj	-1$*+V~�����4���td�鸺�t����1�V��eX�@��^e�t��@1LX̨[~{�O�q���p�0Bw]�����IoojT�B�ғ��B~�?\�\����q�뫔�C�j���'Q�M���1�;x}��w瓹��e/dEռ�T��i��D�W+w�P����µ��־B���,m�^�McEf>ÏG/����� �LjX�@ؓ���	ݚ~���5����74R"��K�ȕ;ǚ�ɞ�һ:�7܀��ܲ����}�h�S������s��ϱ(;��\R��̉Afi7�(������W��(�D�5<����Ss�0����ׅL��е���q�a�����7&�.T�]z�h �p�o�-�j������D,�7��(W�JΟ�c��q�]��*�z${z���؆���DI!Sۀ�䂣��i~f��7
�K�=�}r�����e�9�P�'%�R�Yke�ZvCg&�4.�-�\����������9x�J�e�Y����q@aV� �+!T[�TX�e+ߜ̯}���2K* �����ȟ�UtO�8��ת��T��Z�{Cwé�F�.�zj�b� �y�����G����v��������H��u�-���/B4��|�4|�G���B�+0C����vQ6����ܗe`Wy���2t��?�"���ѫ��,0�|gz*�^��p�D�`r�nJ88���:�` �T�~lu��L�[B�1�D�!ܪ�聽��������3v�R��+~��4��9�;?�3+]&x����
2j@> 
:�~S 9���rC��n�K�q�	#9�S9n��t�XT0Sm7�%��I�i�<�y|��$��H�)��b���Xh�0�ve���cO�a��g��#&5!�6M����k4��Mo[�$E8{7���AӢҏ��3_h��H���s|@��[u��@�����Pj�K�P��Gi�60�}k,�k`�pϮ~{_�����{�7�U!&6��գ�' ^���%'�&������#9`au���Y���$Ǜq����o��4�?'(�L6^�Q�sa���A����3�d��������[�Y�To�,�`׆&���ũ0�2S~����B�=E �{���>�"|����IOh��,om����|x��l.��uG��t�R9S���N��
i
�%�
K<�D�ߡ����RQJϷ�i���3�=Fv���'��?v�̣�Ŭ��y�\��u{�>�(u���l|�+��P`|hݨ9:���mg��E<l��� ��kM�%',%�ׇ�By^r��-L�%���j�dʅ9�?�7���'����qrC=�+)���J���+���N۰@sE�F�/�<�ƗF�[}�����Y��W78e���`��T��-�,��6�&�󺺻 	eKT����U�ކ��N7.t>N�l+*Y��q�1V��$d靰�;���i/k0�����[l^D���C���۠A�gN�_�F�e��Z�h�a��p�T!�e�	��E�D�UF?��&�B5�XPє2
����8�k��?:�@w%{L��W75�@��q��?��w�\ 4��Jǂ�-yU���#����	���\1��"q���d����2-� [Q_cL�2u{[�t�����Dq�$�q$A2�!��vOO�r�gn�L���������5��������cŃR=�F����?��I�ī4�B�c ^��4�A� Ei���>��)�Қ퐖QQ���W0ƷZ�������M������� f�h[b��m%����w�M�k������}zk�8��[I��k���W�c�r�2l@�F�q��w/8v�������X&�`�@���3q'��9ҍ������bV��l��O��oё܈},qP�f�!�H0��\��ߦ-w�Fh�)��Ҩ\��F0�D �g3.3�.F�O{pyp}�	СʈK�#�~Ы˒s���vr9ic���Q�>פ�f+���9�Ԫ����b��br ���<;<C=�a\#�u��|${�5ɽ��B�AM�.��J���+ufz�\�t�u0�~�"�>��<_m�^j�g�2�ؑ�V �V�4�䗒�k���Ȏ�sPjzZ���%P�ގh�
��j�v����{|/�w۩����I���k�ۄ�����e5  .�s?���7�7����L�`�E�E)�I��r��?2򓥥^���.�\�ξp��x��FO����o0~��ܛ��[1��t�#1�Bؑj5 z����V����2.��e��=���i��.��%ߟ�7.@��RN����(E8�.�+&"r�r�zDg��u�Nl$��,�"L�Ƶ�� �i�k/��1�=2฼�T��O��ڃ��%|z�J9���a�K��7�Ζ�f��gh���7�Mí(��|��A.o���8%��u�EMN^#d�ϣ���=:��6ۅ��6;��p�P�n?���G��S��π��6U�9�P�8h�� ����3&ʧ_��lS��c�*�܍��;�]���	���No<8���3�1��l<�_�z����C������A�69�8[�@����HΪEŪ��ӡ��	�_�Ϭ�>u�sg��[�*@w�v?��*�^������E}"�6md\ɓ��=t�^�B:��=S�gvl�#c}-�^1���@�����W�J���jt�Zq��U��f_��s�画#.�l�V��G*���?UC��z0d��ǖb�
���&����w�H���u����pכ�~�o���	�q]�,�麲��f2�T|����.����غs����-���*����������m���U���*i�Ο���LD��T������ƌᬐ>�>�q7Ap�(�A�P�/����5p|9��o]8��eo7����SK`OI�1S(5��v����1��2���1D�4����� �.�}|:�_c�e�_�H7����DS�� ����2�������'����pՅ=�ٷW(y߼,5}�ܴ#l��cӄ������<+��~k�>�w����[���&�F����'3�����	y��`��&�f`�P	0D��?4�]
۸��eV=��uWOψ��4cu��X���~�NeނB��h`����� A��ϩ��j*i���x);�;�G�=��OD=P���uk�{�����Ï�;B� $��n���ҍ�ޖ)���G����o�@-[�A�r�����A�X{=%}����1����ܧ�%~~����3ݞ�B�V@� ��Y9��Z���[��y�#Ȩ����N��Z�4�s�"�n�T,�J���6����| %�3?���3��6$'����[�?29���B;1�&�j�C\�Ř�eu���w	;�6uJW(�}t�Do�`��آ�@}mN�BSq#���h�W��������N���/�\Ɋ���&}�,
J�F�5�-���9e�ۃ�/%%�ڴ����u������r�dM��/��m�ɭ�o�c���N�Ų9���+s+� ��{�Z��e��	)������p�v6��񁘦i{�?�XaIy�||||�!Atӯ *�vR�{Un��Fb�j���%������ /*�@+��Q��An�V&��؟���MT��&��"dk���XE�����{�a��/�����.�Z��TؠS��,ڔUb����ӜN��2�ku�:ES�̗׭5.+jOӕ%+�9,����3O4fOv������n]X�������U�w{���nt2ڬ�9	�0"@X�b��Ւ
~��W����6�!���3��O�ه��v�{�k�8����8�5����:�^99\G~�r㦮����S�2$�W7d�� ?�{�ӈ��?�O�H���5��,��!�*��ھ>*b!�((�t+
�4H��t���) !���]C����C�4CJ�P߽�}�7k�d-�{��g�o�i�,)-��ӄm�6V�Gr��ű�1�\ץ����ˆ��t�	9\.-� |2�����/J��?Q�d�#�����F��%��PJI,]<<&�x��[��-�r�������<��T!)�/M,u���	&Su	�6�QQII	f���6{�Nɉ�ބS!!������WU������9sٙ	K�kT�b�#˻��?{��o���Ԝ�ڌ���2?�
�	U�W������å��=��:�����sLn L�['����c��ʋ�x��"t�W�$CG�1����K�t��d��ڋ�ل��\�c�t�YL򠨐\�G�e�V��� Ҥ7�����T�ׯ_�l�h��#�ֺř��#���w��]c�� ��wV�����b^�xKP�j��pX$�����a	X�-�&{�uttȫ������
�{�U�.��Ω�B.�:W?��� )�U�;�LH�����n������"�D.o,�Ǻ�K��b��x����m�������}�a4r���e�8���Q�3_����#Li�c���=�GA��ʤ�Ä���D������g��8y� T�mVy��A7k�,�h�H�@�\��8��-�O���:%�iJ�KY���?Rz�\R�|�������o���A�F^OO#�?l��l�?'���SW�"�B�����{kj��8?�Қ���>	$K8�0�ak�AW�?T�(���@��
שj��53�<����"�����ic*:�˘h7����5ȌX��tu#��q�g� ��[c�v�kGB�э�+ Ϯ�� `7�m (7dTPR�\ޡeb��t�c���V��m��~�
�j�[�������������/�C|-��F�{0�
hl�B���I7͝�o�J�G���Փ�<�t�:�d���d�C��F���E�W�с3`� ���e"��R��


FM�w����\��&4�{� ������(��	G�9��7Y�L�9X��+�;ou�)Z�g��	��c����b|<P2��f����r��랍]�ȃc�q\2l�����4~PE	�!���[�>���:U�g��ʩU�8��־���yю�N]9�)��%%�bS��B��L�bؖ�O�f6�#�5��]A����  ��_
m%8�?V�Ee�R�K�&s@�_����Zk�b��Y��e���|�� ���%Ă�Ab�Y�k��(��"���z��66#X�.�I�j�D����A�V�t;/]e��jf 2��W�O�X1���g4����BC�?9X�L���_��7�A���;j��}�V��hpQ�,��4���aؘ�����JL�7񦚈W/�|�19��p��W�G��E�se�sE�z/bSJ�I�UrdH5ૻ"�����������!UJK���Y�>��$%�dʒ��!Zsω��Yc!}q�F�&�4�2�i��PI}�G�l�� �)����.W�Gݙa�)�$���U�E<�gv�|�k����x�����k6㷽^�c�,1ZIz@��u�����?���I�(��M�ҍ�q0&XA�|'�9lrA�{A�S�ESf��u�rʞ٦k�����9/(h:$K;���4�v|�Ǧ�� j�n��j�~pϮ�v�Nx(��P�NjǴ����7���dH���ތc���eXD���a���%`>ǈ&g�\�LI�V�\E�N($�}K%�_�ve����/��Y�}�1p�w3䤸(�N��qW��^��j��o�p̌���R�8_�[� ���!\��Y�x6F9��Ny���Ck��ё2mq��m�����0���눿��n�װ�����7&{e[#��}m\!�}|�l|��0��8�ɘ��)߾}�<�oZ�9����Om� `a-�H'���h	��ڰ�w�b[�宅�)T��P<����-6��x���o����pJ�C�S�5u�=Z�1��Y�cS�b)~A��I�lR2Q�t��(L�s�1�n]}x> ��{R#���Nq���_	�N���Iå���-�R� ���@��4�ZmQ���o��]�^���L������gP�	�I�������g�N��4��f�ډ�F�YhK��‿��|aE�5	�W��[�L>-g��1p1v����@���,@:��$�ϡ���i<��N*@����Xn{����WyUb^�%��'�k����T�����w���q�1e.(SӃ��>�V#��m�FX� ����( ��ץ�����k�3���0�l�+y��N��Ǽ!RB���2$yt��&W�cQ�KRv@��P�t婤����d����!��f�q+Y�/�f�j�?�[a�r�|ߢ����e_7��;�Ⱥ�����l���zx��>��c��<�����,���Q��X��x���[�P�f�L�f*�ƈ�Hjo�p�Ou�??�m).�@�ڻ�ʥ9�i�Ke�쉧�,���OKG�oVU	�6��2����@[�9� ��M4�WR1
ݺ��㟔E���䑪�7�&��.��ifw��^sK&؃:�v���F�f��5G��8t�7���$�(d�w�\EBİ��8N��`}�U��&����]�o	�~6�9R�a)�B�1���6@�;���K�\�;h�'D!�ҏS�\�y�Vm\��r� >���N��BY߫��V<��e6,ُ�t���bc�O�]pDiY��Sѥ�`uBL��9s'��z���|�W�Z��dE S-\����`.z7'q���$T�n�������kre�S�C�,���a"��|NmIrc� 7�v���QF�J���+�4�L��~)]ŗ��$;��9�qX��ɤ٢#�r�� 8���$�\Y@�x�� � x�����6�����j�IJ������S)��o��4&؂��;�����-D���,�OF�[x�dd���)4��α��$X� �@<�Dv��,3��V{��nػ�`��V��ɉj�\��s�\ik�r��n�L<��<���NI0���%_���~i�KC�3۸1�ы�����l��Lށ��Y�U��Ԙh����ޤ�tr��&�:'Sg��1�-��Ҝ0�MKή�7��t����d��X_1=����9��[h�a|�MYW	�S"�2Dn/�Ǜ9�2�+��2��ItD�����%�a�9�u����p�I�y3J�0�<��*�.N�|�9i��}��Y{Ԅ�@�yZ��:X�Y��n��e�-�z3*
�fxg�����:��0��	���yq�l����(ꍏ'� �p�$��2�g-�Ӄ[�km��0��$+6��)?�;u��b�"��?+�D��D��K~6y�B�Y��ȑ�W���cW�pm�`��>c�A��7EQ����-���f�����$��6Q�`
�� �H;y23(by�RLǈ}M�}����4%b��O�N͙E9��e#�%N>�e25`!a�Y��[��x���:�b
���5܍��|��=�"�[!^��{$�����	���zҨ�W���#����wR��(�X6mֲU�����{����~�P�1�r��{�����I$P�(�8���n@����2���9���T��O� s�m7���Erp������Bӈ�ΰ�&e��!�C �m�R�%��7'�Ʋ!T,k���v� �3�¤����ӏ<jLآ�[.�o�A~M��	�0R��8x�&� �f�P�k,��Ǖ~�X+��(�x�w��j�2�,{ӊ/����	�]�O�<��fШV�i Ɨj^0Z�5��a!�w�"��G]j�������O���BT�z;
�R�;8dU%����ZX�KBG�b��
�ȭ&�s���|��;D�櫤�/:�R.`��oQ��"
 h��>/3���~[_qg��Lz���E6pYI��(��$���kvF]R���=�!
�Y�uhΧ�����ۧF�8�C=u�S��Aۙ��)�~ݒ�3jW�γ�"箸�.����թM��l'���dn$�A�6�7��x�,��ߔx�c�Wn�esJǆ�q�Q�U84k�)0�����5�z��xy٢� u�&yו
�O:/�U2����)4\�Q:A�qJ�����
%c�$lt��<�v��
Q�{�����sBJ�._���N1�ϙL}��|�S�{Kv�K�O��;o��L�S��ce�W�v=�*�WZ�x���0�e�����u/���]ƍgf3Tl��q��JГ"������ |+�J�����G=�D�J��]Ж����rQ�N���Ǫ�1��\"?�2�۷s5����`�(���C�<\�s����Gtk�G6W	��S�މ��/1^�zn�T�9{�OJ�; ��播�����[%;�J~%�H�������_�8�?���O/[���/Č���};����yd;Dݺ|m�V��s_}Q/ J�$o���FL����v�u��Hߦ�6=��͞xr�q�i�%��^w���qg-� *�J��#m�R��
]�RZm5/u��ƍa�"��\�69��so �v��-�z#���FCArb���ˡ�A2�u�v�Y�lʫ)��q��.��t\jH(��9��B��̒��Fp!�ʗ��>���y�)i�IՉ�=�J�(jW�<k��y�x~�C�A o�#FUS�i���H�w&[m%^Otp: )1���=6(yS��>�SO�*4�f;v�Xa<�
�j%wu  (|����!�/�mY��av�b��-4���a�E?��	�3�V 3�+|s=���o��S����8�y>��u��?��'2�+��;?c0����>�*�ǝo��M���$4-1�_�e�·���W��c"ް�*4�5�Ù��x*>�F�x���C�?�9�c�k �|�2��s�t���-^_3U���"������`K��'Y1Sr�󛞌�7ӒΩ���a��-$���T<�'C�Y,7uH{Ow(Z}%���L��u���d��s%�%���k�7/��ci4M���C�&?��k�D�V�}"�'�^Ae,b|�n��o���;p_>8:�\$��d�H�Bߐ��Ҝ/�=unD���V9�x��qu<.���l0��/!��TQN���*�Tn�#�ψ#d-aɜ(�N�K���N	�~|�����*R<"�N�OW�q�~s1/�\���(f�qX�&��X�=���O��ݝ��K�"'.�K���G��7wt�Cm��u�ׄvl��YXXX��7����nQ`y�$�05���� �ɑ��:��U�䱙Gl^������5�d�X�7�V�&�3 �uW�b/�^�6J�G��.Jp��G�cL��@<ϴ��o�ב{��S���ף}���U�M�����zg.u%��=�f ĩV�Q";T�12."T�o.k|���Kc-�"ԭ=0���*"�!G��+�ǯxx�K�^{�e�k{$�8~=������������ܕ��)K�&�z��+o�\(�}���,��S3灁�A�޼���8��jc����j�3λ���3� G���9�]21Ͳ�KpX���E� �q�:��Lҿ!:a�>.ǠDB��1.�aP yv����ʀ�y�~l�]f���������O������`uJ��f��^���˻	�/O"��}��ƻ�Qi��V�ջ�.�68{�%�8��-*�"+�\�,+:`�vS���8�dN�(ބIv�)LI��9���'^���~����@�� �Аgs��t{N��x�{�U�]��5_@�����f�$��E������R�z�-��Q���֥�ƺ�f�;�Ā�In�B=W�#͛��rpm�����ȇ'�dp�Ro��5�v��z�P�5G<��^|a6�W��׺�~���E>�Y4��1U� p��VeU�bY6���
��to��iU��
��s�����@_�9�I�9!LE�$)ve>��&v����˨���p*	�$�� ��x-�n+�@��݊���Y�Vx����/���}��Q�'nO�l�7��jG.�h�)?5��V"��ƣ�|2�x�����_p�N�ȓ���ol���~�3Q�#�2yp���:CN�% EN����7E&��+��f�fP�r�Y�+���_��"C.��T�T�+̡�/?�2�Bk���S�פ��pr�h�:6y�ytt����H�����eء����D�ź*�3��_%�+!����4�aA�o�&�
c}<x~q�qP��p���}�/�~YfbTi�m���~���qR���,ߵ.n�����[��ѱD�]4��)�ٞ<N()Y�[i�yc�P,#�k���C��cr�nI��� Z�*�N�C���;ȡ+�緈ZZ�UY֜���
��!\�R�����P���.cS�~?*0Vn2��_9�LDp3��'��H�QGw����7�H�6���)|���7L��ll45�mqQ)��gdy(��H��N�Fp���&�R��!�7$n��H@��X�L�S֔���!7�Oo������!�?�o�o�c3�������d��3����a��`?}���e��>�=66x���H�p�?{�HK�����l��������Љ�ZX8�{̢�U�������S33���gQp��d�G��z�ផ�ryv�#�z|�OP�^'�s��o��;m{ݘS��.c8���ɢ'��mć0��hNB,��U2��*^!W�d����):U��ED�,!h��}��.ԡFZ��T#�ñݏRV��L��u�Y�yëJr8cZ�V�e�45���B���*��S�9wc�L����"a4թ�t����p:������5;#�߽".�|qw�UZ#�&iYvS�.����l)m{��Y������_�b�^Φ.�L��r꾃�ѿtΊ���]�R%ا�CGO�)�姨+�)+g�uFа��`��m��Lq8�w#��I$b��Չ;%���+�{ꃛF�w�a���J�����/����X��Ka�������R�11��'t#���(g��� ����?+�b�D��������/��#Ww�ɞ��1}ݯ����@q�֚0��L��oI���N���EF�U���b��l�b{��zm�!d�w�Y9��Q�*��09���턜�z���?��e���Ӱ�{�x��w�f�7��l�ě\5�n\*e��\�VC=t�ed|drA?-S |ٰT42�@��7������|�ω���2Fv�d�uL�捂�g��dvaAd��G�.}�l`��+	���vi5=�5½|���B�է,m��td����^�%�/S�ꨕ�w�%�u�@Q9�D��@^�Y�N�)��x&{��Ң�U6�1��}�3Ipd$^�5�Ϊeo�1��h5���INJJJh9Zi!��s����;��]�p�4"v��<@���[����z+�8auf�.���j�9�;ZK��Iy�^5�c��t7�zh3��;� 2U�+���}꣐��=�;�б�,���)7F���j|�H�Q�q��\�̾b�y0dҺ��h����}|�$�`,������b/���(���(��4�Yr>���'טkvK��+gn���ǝSN]�h����^Y����.�q˗G��\�$%%�^���p$��TY��5���_�GY6��X�<=���{���O"�� �51����lш���r��7jrI� d4�x2�FX�Iq�[��$}�)L��x~+��,�o��Q�O�t(���������`��Y�϶�t����m|�9'&�4��Th�3�g6�
�z�br��*g,!6������^y�=��c�/XU�kh�sc�cYZ^��{��#z%G��.���ԓ�Dn��zG'ώ�*�8�]�4��B�=��jF�o�6���EqL��,���\�OINV%,|Nd�b�;���D��R��i�A�֭Ӵ�x�)~m��k
8������J�~��������G�2þg�v�.�s�J�jp?��־dЬ�3��ͷ/PX�2��wٹ�t&��o�4�A�#$k�F�)(�W�Ŧ�t��Wl�;Hֿu\�����v,�Ȅ�Z�ڐ���Ͻ��������w��(]��#	a�΢9��nL�g�,O�R
�U~��^|k�^Y����wcvn��Z����Z���R�V��q�ꧬ|�?Ku���zz��1�}��`?e�|��:NK���N�gAX�cwm�_�jNmQ�"9�i��z<���,3>�鯬98��"9��;8�x���ĕ3H�۟^���XASM�*6z�;ȍD<���&ώ.��v�K�F|6���nF1�C�A�}�A�+���7�p����T��UIX�6��.Q��.��a�g����r8��.+��nR�1�t��F|J*ۻ�sq��1<c�L"lW���PW��677ˬ�:�"F)� +�&��P��4E��k�+��u�J�$#T���U�K24�e cQ�v���U�]��7����!��Rj���� R����P�9P:GM����Ɨ�}	]�,V�2<����V[�g'7�6�7�j��ؗ�g�1�+:�H�v��+&!�L�~����=�ͤ�Q�r��g̗��j��������E9n��Z�P����8!���=��t4�_^u���"��TK�iU)ZsPB��d�@	�$�\F�KX��f[�"?�S�阱����T��:�3��z��|أ��	�h�������m�+���y@Ġ�Ln�%�����YP[[�U�&'�
��}Bdu���n�V�tj�XʥU��h��6d���,���8�u��Yz��Nu%�9,��cϢ�v�P�<�]�;3�6K��?�N�O���G=_!�6"o
S?�:B�Y��K��qq�0BR���c�� '��ӳ"�$��R� ��N��HKZ5L�K)!v,��J:�K�V5����*d�.�ua�8��|���CC-���B��������
��-� &wY��*\ǳE��~o"��ǰvw���O����w�k�g�-Kv��&9p�]���&����:�f�]Ч\��v\0����⋩�I�1��Մboԝ����ۋ�A�f�>Mɟ��1��GDFf$8P.��6V=Rj �?�fv{�*��7E�S��7<�>���%���I�_;�����-��@&Ջ����՚��V���a��O����6qo���Xq�ԫ�RW�|8Z��e~�NBpP�T���	#?�������e*��������TJ�Nv
S+ ��a�4�*�=��촯�l�Y� [�4��j|�/x�r��_:���ȸ}ÿ$�lѧ%�^� &���pS�G�t!Ŕ��C����@�B���A}1"��-+�g���Jpx���jOA�\�/]�|X|Z5L}p�.�|>v�H�O��X���	����ş�C��hT�j��0~���m[QG3:�g��k���N�V�wV�H;Q�^�X�ˡ-��O2YM�o"�ꁦ��07����S�B*ji�T%#��(���roDڬ���侫�A����8|qqdv�a����H��%1F�B���J_�Q��L���Ys����T^/��y��-�)�
�qy��2�S�%u�k2J0�����$�pO�6��sd���N��Y�!8hҺJ�����hE/X7���T������D�W.@�B;��&~��/kB$�,ȃ���mN!Cp����bӱw����]�
�L0J�b�uR�+����-�t�����u��"a3&�˝�"�2�1����uUn�1���-�!|U�[(�-�L܃/x���w����?�Yes��
��_�d�q�h�ڳ�q���e͓�<i3r���.��k�;W�_5F�����\�w�^�`�}�qE��,�R-՗����g�ǵ�X��J<%g�+�^�l��oVОx�����N�}����4�h�Z
�D�mo��ֳ��k�0q$厖����䢪D�&|�*=$����$�U[�|����n�Y��nv�i?N,&���R٢-n=Zì'y� ~:���$�ls�n��PA�����@�]�� �~�@xK
��r�6���褴�B�>�Sԍ������W$���$Q�m�O����B��%	��9�T\�3{�5;ē�bj�u�8TR�K���o�a��U��S���G�Ʀ �w�@ހ����c	���o�&��,����ܭE�LI�K}�x�x|����I�OIc�Wʫ�YUޘ]-��M�T-��-�r�Y6�����x}�+��dn�:>eo?� �E�ʸ9��*p����T���PX�����ܣ�=��	�j��l³G��c�uEȪ�|�����}{���o���@o�SiơvFm4k��jO�OO�c^:�D0�e477g�!��q���K)�Ԏm��My��j:��l��h�5��f�k&tN�|Vf�$�V��nǠ��ѓS-�՞[�褣��`_M9{� ���
`l0�f�����d���9>�2��$E^��s,�l1�?B5}UZ�\�^b��>��[����k�;���u�4��3�sϤ���>aau;q6��ck��V�E��W:l�e��X���ly}�T �I���G Ϩ��|�`o��a���W^�q=a1���O����8,�2�7o�X�:��+R[NR�v��ұ��Q{���a�&�Xl
��_&�Y�I���ٙ)a��yi3�`�Tp�ʠI�u���r�ol��(�,\��d���*F��v��d&���a4V�q��EA���A�h�i��ā���
w�������F���D%C�n< ��)���y�\$�P��^X���
8�x���>.{�	��ìS�V6[z\��X.�R��Q����)q�r�놃. 'R���֭�H��K�#���ꂂqC~�D��]��`r�#۱ҍ�Ý��5|����S�e�F%Tg&�$)X�:���fj���M���Ig�8��d��� K,�.uĵ�oU���k]c~������2)�f;بx�;^s3�,,�˴��3ȳ^��`c��qYC ��Q��֋{	8*Nf���wm�.�� ӑ�Z�hw��`K�/�37��d�"g{1+����ͪ�j�p����g�<C���}��\ER��5�+l�;�z��0�׈3�e�\�8UK Cs�Tj��S����-I3W�N��o޳6Lw߭��n��ݕa��_�6)���;g���b���)���l�B��\�B��_~���v�b
6��{��jI��`��r��$��@6Lf×G�Sؓ�3�ձ�v��qyvR�V
�*�ļʹl2}a�/C:gTB�ʳ���TM�<�z9R5�إh)��FM������@#%&�W?)��T��J@�&��x��6���k�7��`���t?*����N���� �,$-Rӕ�x�Y�7擔6b'	QQ���q��ޤ[��+J�f�>�LMJ��7�������+G	
 n�YEg8���j4D$�ҪǼC²�3A͆���uX��1�,�V`g��Sg��P�|	�E A@�[�5���a$�����Sžj�7r��[H�$�v����
XE���m7w��� ;N�֕xq"!��܆�z����Ϫ5#y�����4���� �G����2�ֺ���JO�j��"L����|���½��ŝջ#.E
����0 ���\��j�>4�@*��y��g:>'���d�W��m{�w�s�ԛl|���H�u��<�9`ᴕ�ZӾ�HT����aJ��vNbib��(� 	"�߄s�l��� �c�Y���闳�L�;�(��f�(T*l8q�x��g`���LT��\�!�׻��+((��D�A��^�����))��-��о��7��E�:7�;���P�7d7�ش��������^m`M��L.��`
�UGc�.?[��HU�'|���J�7^����C

H�[�Ei�
c�t�Q�*��(*�嫼������f\�����&B,փ?�7<rr���|��4�̶s�yI��0'���0!q��[˱Y%q�wW"�բ�a�!�BL.��^R�!��x����7
l_I�)7ۓ ��{,�ux��Uk�1��t�x3*']G�P���S%"}gy06�
�
p���<����FO�.G��������>4���I�w���ci/�E����07�p<��[�I���=1� Z^n��Vs���+�,7L~<�k�9�<���E�"�d43�4���q���W�Q�^����޵;2�ٰ%ʱLv
d����DC���s LC���
5�p̷���k�y>�{�n.ݯ��k�<�y}3�|����g���t��R����҅������MVɂ>��2��EAuV��}�.Q�2��\}�@��b�$ ao�e�@b1�o�G�F�����2s�=�qMB@�⫹<%�}{����]�^�D����[�@� %�4B��C;XH��o�WK��vE�n�"���dŤo�G�؍�鏗��d�c�Z�jHٱ@��'���GgRWt�W���=��O���9D(i��ٰ�J��h��w25�){���KFdu����_���	���Z:u�e�3�����ܒj�lT�7)D٨FvZ�[�x3�W�c�Dh�R��x|��r}����;���^�RI�jZ��������~B���v���Y�����&��{7�c�T�����|����w~C�5yR��T��M�]�\O�+�S����������žTY���˙ ��6������$0\8�#�t�y~��㞠�3�f�NDw	�t<���Tc�:B3�2�on!�}���H-�9>�� �-4S���X9	9�I��0ޜmW��J''�ZS��,��|��q�!��� ���ޘuP&����I�5����Xs5O��~�nd*c����8e��S���w�ư�k~�n!`ܳk��v��<�#�4�v}"?[.sɏ*!x�<hi��`�H M�(ߘk")T)�o�/}����&ù�����zU���^��o�Y��#�F�F��O2��=`���*�_ʛ��]�<&'��;j��. jS��C�tz�����t�h�6�a��/k�t�,�U�Ӹ�D����$]\�N��m���oV�眒�ⰰ���AFi��JCkP�f�7 ߞ}q1�� �T�յ޼�`>���|o����`Ô��$[����8ظw��1��
ߣ�&�/k�_�Ҕ�C
��Ў�R[k)�[�	�Ր�I����X�И�6���<�}�w,#�;�q��z���T����vG�
�T"���D�����6��j��<�"���hP����k����^=���;XS�0�o3�Ϸgҭ}��NA�P�{��r��������?Ȁn���5���PV���x$YbO�����c����
��ޤW�̬ 2��u+'7�%�
�S~��/����71Q Ji��Q�g�}�?X9�
v�=x��v�I�Y1lz���ai#�3\�V椅"��i�Bخz�(�)+H���$[tm�u����.}��h��7xO:r��e�m���rNK���SJ�eED��-�YkDB'��0�����v��z^�o+))Vxd�	 }��u����*�݇6[]]E�;^@�Y����1�^&��D 4�1�UC�t�[�SԬ�~շ������&�rO8�Y��?���צ��ԡ��,|{�O���?4^U�����fQ��e=�X���,w��:�zpU�����#�_m���N(d��Q�*l�)��L>�w7*$$��P�uf�d,eä�5G��qq�) k����=`s\���x	>ܿ2\��]��h�s��|��F�t"_+3 y���*���c.�	�V���u$��&zYjǣy�=�г ��|^��ǝT"�{�-\�b[����H$ *�777��qڮD�W���'�u6���>�լ96e�6$_h����߿����Lk�dd�*c@��X�y�nݺ�8�MD^QQ�^��h,iﬦ��N���,�G��v��8�AB�RJ��Ʌc�Ō��<�T�}X]��u��jfHDkC6���hU[�+K7@�@��i��dd��6sݿ�^(---d!��dW�[�4[�Ϯ���'9c�ӓC@.���˫������{�,'���fA�k�N�a������Հ�)�n����{L���`'9s��ԏώ�;� ǯ�[�E3�s8o�ˤ�_��r�9�Rб���!�kT<x�d�_�-�	v?(��$B���c�,���`[Yx�i�s-�>��H��B�c��'�<g��,`pD����$5ł��'Ǉ˭��B'�;o��m��� /1����e�05u�6�U\~|�@���K�U�S��a>����s��"-բ�Vl�Řu;�m����6�y�j�ބS�ˡm*�t����rVf��Xvvv+��P� <C2tr�#�J�� 8S ��vNN�a�=}��ꨒx���bD1�G�b8-SFFF��	8'��m38���5�M\�u�73
G�å��SR��<161a�����Ύ����?��Ossr`�v4Am:�>  �u�L<i7|+��mo��.�]"�~e�J�;=';�Eĕ���4�"�Ѱ��.}��Ԥ*L�S���S߻��K�r!��!� �R�.���L����1�F!����צ�� K�Ml*12|�E8����\2�Z�n��U����R�����k��E!�������>@��� �gȍVGʅK���v�� ��B}�gJF0��T�I��8l5��/(��ʋM�N<�E��/�!d��㫝�YN)����C�����G�������#����|H�EP�n��O�t� �y�r���w���G������~�ip����)cO_�7a��p@�G�n��H�zhՖw�W�dt��1�m�}*�z-�л�oٮ�0��W��R�}뢼�-:c`�4HI�߹ ݏ�S�X�}� �X�~w �LIX||�l��.�3�-�[2�тg�d�ƕ���v���Y?6�B�da�!��tTk �e��^�[e����}`�*�����<K��kԩ����n����j*�8�zxu
�1����w���\�O3T>|@S�D/	���b��v{�J���_<Z��ݻ���SIu=F=����<o`L�����h�7<f�û�s}�����ܫ������d�M�/p��ڱ�����������A|D�T��:�(��KE%����c��p�l�zhR��{�
�n@o�@_�����-e�
��5;����H�8Ȓ�A|��%_����.�+4/���{�V�����5��&�;�Ik_�K�޺����A����~��eٴ��x4�t�k�b#Bm�������f��,�?g�l��꠶��,.�<�%�6��_t���o���$*+�/�"W@8���XG!Wт?Tf'i 5	+�p��,Л��Zz�� �#�,7e���'1�/	�K4���\���/�%^� J����4-~
�a��$�J]��K���)�/B�j���a�2Ia��J3]l���v|���E��n	���
�65gT��R�n���YA�X�&gk[�aU��v�lBXX��S��#�޻�8ᴎ����o^���g�DoU	D]&"C+���+�X�Q쪲|X:6���͘@t�V�4n֚��%ͅh�6�t�m���"͐��sa�tc��5�,��|~�Z$g���9�`���]j���5l�+̂��u�`�2�[�ט������8.�Yl��t�)��w�1��j^�b_�ÂJ.<L3�0���Q�������D�;H�V�(�=3�k���4���g�@�Ʈ}r�p���7��:`;eն$���B�S�!����n��!��a�X1r	#��v�4"�?�&s�4�j�꠆&������-�?���_6,gV(Wm�R+q�S')���+'r�L���� �*�[��%yYV��i�J�o��@�z.�w�9?�p��_UG��Wp�;P:�M!�)b�J#��~-�4;�-����*�/~:��k�e���*Jp3|%��sf������V��g!��	���F�QI'�-��F�ᕓ�j 
fP�?s)��aq�F��_Z�Ӎ�T����'<t��u�+jʖ?�ֺ�[]󕎐��<0��<�歾�X��i��\�f��3�xO�ioQfߞ��0���	9���#9�o��e�u�Kw��)6_��UسY��u��d[	�� ��j�H�ؽ��a�h�C��z�Mc��0��=��.N�gV��* �@��kT�3��=0.J)y{��'��F�r�6VUM-`��e�fi�������*1��4��G�1r�Hǲj0[����"t�T��۔�𹂎��r�Ɂ������p���_�X��y&g�0"����C��c?#9��]\�1.���>-x�59���l���ݒ�+�#Y���7g�v�f7�%D���|9��&�ͳ�=W��ښr;��X3f%:;[ҥz���ڗ ���H}�Rk�E��r�����98��Vm�+F����ҁ�(]��R�W��R�(���E�6azc[�&�=����@v{Ip-��!��!@N�h$�UW^��oJ�V�6�,g���y4&�����>�	#9C�"��b�D���=B���(��&�3�����ǝh������m�ćP0�[,�s�4N��|>Ȍ����HwY ��<ŕf*��r]�I�4�ˡ�x�a�~�	F����r>������"Ξ�ѵ�e�F�Zn��D�;0m-|���eg&�����A�kv�����1Wi/�������}�^�*K�Q�U��H�a��C�%5�Jok)��ֵ�;�=O�:8?�1��26�\n��3FRJD%�����B(�FW=�j[��B�� )ɨ`dd�w���\>XH� tٲ�݀O)�^4����(ۓ�^��8��<�=�<Ӹ,#W�s���A�8Z@�ى�� �Uת�v������3��'<��'�����TUc�N� pPH�"5]ă�~�����Z��0�x��F�����Vs9yeZ��#=9�y[dz�s�vHZ�7b@,�0�Zo�GF��U�o�Ef���>`ym+��[&��B'IVLd�Y��g���L�9��u<G� V(c�-��U"8'�E����I�/�����&������,_�=R�!S���@�ՅG����9	�䨖gת���eW����4ߖz���X�
%0�o¤�
�6&&�F�T۶�ɵ�?+��GL�a��e���O}� ��L��ϟ?�iy����������a���j��:S�rT�k_�ٿ�X?TMp�"&$�O޺��@Z�I�B��u÷W}�m;3J�� �Tb��qr�o�o���C%o�/�#�!�T�vt�,��	����[ 2BR��w�� w�!�S���=��-��x�MO!���*�A-��"��X�����g�r����KbqHa�ƚN��Af���*�Fdy�Ob�����͹�p ��W5B¢p11ج�%���zݽ�(����M���i�� ��EdL[���>�LB�9���Q21tɣ������?�)�����"+#�C���#[B���J���$+�d�B��Ce{��{��p���������Ox�_㺞����%L2{���Q+�/oe{������g��%:�I��>_�/�2-/.�J��D��}A�P�@��-�
DB�9/N�n.�&jpW��A�����z�B��5��@dٴ��.g&����YW���O���:�k2Mۣb�k�O�]&?C���|⽤�m>+$����s�F��"����S*-��>+�+qH�;pܠX��G�=a�`��H��}ҍ�"z�Ϗ�������|�d�����3ƚ��΂i\�����������	��w�*�����"�O}��ج|���Vg��5r������T��;�����ȉk�`�3]�~hbz�wu{g~=ñ��JN��N�Z�!����o����� ��������=�!�-�z��x71����aULX��,�ӗY��Z:�im�n'��Y ���"`�4;;�M���b�kHYYY^��#����,Gj2Ra�p{o��:���jl�(�/��Gq�'�}�l=R�a>��ʌ���)�8���o`� ��x>��3�juk?<��<#��8�a�50{����vk�bY4�@a���`P��~_�*;�[`W�]nCxs;��X�x�va_�c>ctz@�-����:[�w�0�2��00��H*ݲ���bJ&�&�*S�V�4 V~Na�o����\� C���\��/�����a�2�ĕ��� �*�7GQ�J�"�:��������E�1�ʅ�u��W�[t3欏dv���j�х��=Jh[����վ3���p
�E+x�<װ�@����&�,�>�����<�*�9`n��� ��-AA-A�s8�U�ik���%Fz��q�b���[;���J0�����7�p���������4`�tB ��Q�A���@���Y�O7�/߇6� י���=�I��f�ǼD<lſ<}�8��tU`Xϡ��3��UJJ�3�ev�qx}�y��~@�"�[C�WW���� ev�4=p�Xe�N�bh�~b��G�s:z�B�,S��b�9m�Tm�r-���z�%�x�=F;E@��O�zb��V�+����s ���ϣ�P`$���\LFJ?�H<��`�ң QXBs�Lz�E����}��!����q���ϝ�����,�l`�qz�q=���qH�Bp�;W͒��F���t^t�-?Yo��0��XD�^�N�,�f#C}[�L���ɭ0�o�V~��<�<��a�y�� vWvN�c�מ�C�Ik&ֈ���`�VIÜ?O ���l����{���D!��P�)�=��	�v�SC֚(�b���ᮉ�9�5����&��Mb[��������P�̂�Lz��AM�B&��/87!>�=�� 9�y�5;��|o]��7��5���"Y9_:T�8!���LA��� E�(� ���C0�����	�i�Q<�>qY|������V�����$�2��u�q�@$֦��	t�-g+�_%�h}A���̑�8n^����d��硸J�r,D���P��ù���fg��?th�����KM���Do؋�)�0��6Ő���5��y�B���~-r����:�Ϋ�N�6���T$���R)G��v���d���S5BW�q�1'�ө�����w+��,�wi�î����'�b�+��lzlF�$M.��K����e�����_g}���Fύ�B)��
!��Y�<�ߒ��
?؅o���A	�/���l�|�[�"��W*Q���
/d2��;1U��Yέ�]�=M�f����#�Qz&"��[��17$BZ�ʲ���r��BG6è{����t����"ց��xڄ����՟Յ�
��^�\���g3��-�i)��"��.N�!�g�9������vW�Ӕ"���_� l��������XJh�4��-s\�K��z����4M��Ϲ]����Jo��*�ś�
(2R�����<�%
#d����]����뼪)�oF���+���zR���OK�CI�����j\��~h�p"I�^��jio[���sM댋l�k<����e�=˸����鄪�:;�No�W���s��m�#ƃ��Yj3J�)�����dHl��z�u�Z�3h8�7 ����8��=L��
	��Z?��5�鱈/U�w~cK�R%%f��8u%w���:�.7�����UN�z�+�r����-6�Sn���0�R:{CJ���1�p���2�z�����I=R�H����Gr+�S��aO'w����ON�cS�΀�o���N�l�_��t��e�~��+�&ë��:�L��>Y�)��/�|�d}�M9�D>X���M\#F�i�hY齡,Ów��ev��]4��'oEۖA�{��cA�VV|�ǩ[��g{_GI���*v����Y��M�1W�[���Υ3�=���2�f"Vx՜��\���� C�1xsd$����������M�[2&Bme���P�ld� )�r���C��s�o~@�@j}�����q 1�Ǽ��0�_�r�(ի;�0��g��N+��$B���L��|j �T�˿Q�ѺҀ���S�{�lٟ��+���jc��"9��'�H���^�a8�M����ٹ9�Y1��߽�S3�̌��5Uݻ
*rCW�ߚK������?L���x?j"�!sG�c�uGw�2����w�e�V�b��|fJq$RǏ�˘�<b.��l�\�,/��_g��S��zU)�������Z�ܷgY�+�x��G@C���I;�$�3Y�Z��ڨ�a�5B���D�'Ӿ�癶ju<û�J�:h����`�*7�\�~ޱ��������PV[�w�'Y�w�v���J���;���g _�<�3�8zp����mKz��/��ٝf>�,~�ok�i�R�{dᖓ.6*�G�oEp���cޝ�)	Ģ���T���TB�L_΅�_־�u�(I����-�^�+qn�$�hVi���cd�7R�#��[���'=��ai�b�%�U��~����(�3��hͳ�ҔO��`)"�Σ(3О�S�WįH@��Cȝ��jdl[܌�������]�3�������M<�~�b��OT��w0�\�B6"v��T'�IOV�Mm~/u�a������m"=���Ԩ�Q���d�D�R@~�ku�:��?�xN(ׁ�,��ғ|v�m~�F�5`O*��uKƤ ��l(x�P�V]W7Cg�˃�ub.] ���"w�y�Z���fTAEҮ�ˁڪh(��h*���e��S[M��T��l�i�u�\T���5-.K�-�:36������8	�t���w@�� �}JW��9��SV�r&�a��ye���n�WIz���v��S|�N3 c
G/<uSz��B�ҁ(�|��IA��ʚM��a���z7M��#;-���V�r�[�D�����A{Oׅ�,��j��h��Vn�t*q�ׁ��cn�KٺA(Z_�`;/�~^�����������W�b�~��ZjwO��W�+�bq�B��L����&V�Va�Ǔ�We�J���3~8�Q?��x	ߵ�����7>(qj[���d�,v_~9}�τ]~�D�0�v�ѕP�n�l����/�G�ϖ^�r�aC�#�:��ٞ�E��?bDu��l8:���$�f��-!�s�,�����aBtt;8;;�y�(�n���$9����������k��u���!wk��4w�$ux�R�0��C��4K��%��c�%���Ș,���/D�|����dO�#��y��+H2�W,�e��B�W�36����Q��F ���[����b̮�sC ���мN���e"r��Q���WT��ԙ�z3�����L?��ˬ��_���1-�Ztʺ1�f�5�����GL���#���<6���C<N�]j�P��)�G3ї��2�� ˬd&����zL��NOtm����;�;�X�}�g���j�E�ZTO��ﲔsB��ܔ����?�B�8��#�h:Pq����b	햳��ۜ-���m�huo�v�ie�wX(*y�e&`G��w��&Rr,�0R��`�����L��:��v��s�@��k 8�:88(?;I����f���u�����  9�n�&�1�d�����^v��D6��M}�%�&;G��)[��2�z��z-S*�	n^u�RȎ��"��@22���	� ���)'���Lh� 11��45� �j�,�93?ϟx��o-`�1`�~}L�FJF���DL��Y�%=�ff[���-���F����N����r�6�yxW<,�z�J�:��T:|�V�M wblX���\K ��T|��p�4J]	`���7����݆�����DFD ���ӯ����W�H�ae �ee^ �\h�km�1�ѕ��/n����K�9x�o��x�%��
�񥮭c�9����Aw�Z�$�N��l~�TQ��Ȕ��@oW�|��/<��a�H÷��%ϊ1U�mjRq�z-THc�{#,f��JJJ<�
Znz���HU8e2<]�C/��͈`��K=O�OzN��R��.����U$0dc=��lN�:��={&?5b?�bt�v���W� �Q;�7�����?�q�_�b�6��@�o��z��Ib�e��U����(��]����
�u�������*�Z:��"q� � �9���TO�8��Y��Xʷ3%N?o�GJ��Dw�n!
P�څ�7@]t��T�(K��ΰ��(yæ^F����?t���}��5{�
=[���\2P,;�v�r���z����N�Y9����ɓ�!�y�ZCKk6�ed�~�1g �e[�m�elY%,������[�;���.4�6:�p��!���w M���=���;4��"o
�s���-'uT��?&q��9(�Z�?�䕏9cR��g�Ie��֚����AZ�{��c�1|�kYl�Y��8|*���D��ї{���y������9�Od�nӼ���dX�����5i`c��&8,�`lS!+�-���b28̼"-�w	�H��o�.j+��`�*('X��L��u�������3���0�@Rf)=�M�����^rQ�9t�[B��X��!r���ϽC�7�31{� ����{�n'�\b���L�y�.�����T�*�f-֟}��'��];b�ya�#�=���yQȚo��y����**)$�O�]�*�펏��%��m�J��ws1�	aY���fE�����h��q�����X��L��.�s
�x�h�(�W��,����~��aǅ�\`����V�9���S� �w!�*霿��p,��JV��O`/���.��O�o�C*�y��w$ͨ�\|5��&��~h�)�Ce�[�c@,�q떲��ّ �t&{{�xl�g��8��͊^� 9��f�x9�y^��4g;�%�% ��S2} OEYݩ�Y�L�g�]Y{��7g�sF;��[Zx1����ފ���gB�gvf�a��V1�����Mp�+6�AU5�/���"�3�fm��(!;��&^�,��Z���f�K�����������A���6�5� jd�z�T��K�d��B��)��!x;��j��.�ٱ��8+��bCy�'�P����ٝ�S�U���aΪ�K�	-��q)KD'/�� �D�� 
��\�g��G����Ml\�)׼���������� .B-@y�A��?�V�.V7F"U�)��F�0F�ʘ��ˈ�Tl'���V���D�,W�T��
�ǀz�H��)�I=�I���.>�'ru.�:�˪��W����r�y#����d���w�B��X���	>?6 ����U���Gd��і���)6�`	+�T�[Ұm���,�n���墓����h�u���Di��}�������E�h���T}����آ=�<i5 �����r�"n 	QF<OD�Xe� q�t���ۡ�^�̀��>��q�����ωS5��ru@Lk
2br_
��q��	hO���0b�I	ߢ�z��U��##�L"��Y�Z�y�ށx���o�{#O��j�1'��p�b4PVY��C g����Eh����wS�R R{8�Y�)����s.�w`S�~��r�l\�I(�uQ�����=��*���S~ĉ�d��]9�},ਗ��|j�?��2oe�y��W2jkG��׿��jI쟋4j��Ѷ�l�f��<�rL�}�c'A��k�*=i���Zg����1�c��Et�B�xGcm�����_�z>�����X��P���;0`!B�؄�VꚚ�p`�}���E��*���*�uB2���Gm<H&��a瘝de{#8*T ���">��zWbs��`�z�JWR���E%Kp�'�{FQ���3�r9���_���)\8 �tr�,�?m�8X�D����-c�Ȝ �F��Rd�4�y3�3J�	��@`ݕoed�1���*�dK~6}�5�Im�>��3�%�����s�F�5q�wh�}����g�<�*++��6m�4�I��ϐaUL��K/����u�iSm�^�NK��Uj���Y�~���pҀ�v�1B�Uu%�v�r}�cH�Q��@�K ����/Nk!ߌ<�nQ�KJ1Y��@g�982a�'B�Tn1&>3~�E�{���V"�jڍ!Z���IO6w���)8$w�)��9e���T�:��	Ł  �wfx��'m��H�x�;ʴ���b�t����)3�[L��b/��,,�<R�����f��`%:��`wB++E�����e����«��x�퉒ף'F�דn��_r��7,;W��R��I���9�p�RK�UU��I*}�+,���3�t�f���J\�o�����}��p�
�a�,��yW�����w�=q�Ny��+�������v^w1�!}b"q�����%Zú.�5�����NCA%6��U�/v��E�����'4����;(ȕb�?�Qc��/_L���V�`D��n�r0�� �����m��,ws,����`��R���ի�����e�U�����y���̠�i�����>���V�r��/:��aVB� r:_(8����8�y`@�BZ֛(��/�m����xxT�o��pLzo�g�����̨F7f�NFX���7�����g��-ʰ9����h�v3?��z���|�`���	ۄ��(�ͬo)�}~��ou�d�	*n���_=�<��1��y3��W�c����@�4J���k�?�㯜�Α���>��6P`Qd9hp��*�A�w&�ܠHb'����RZE��S��j�O�*�����pv��sX�y�8o��Eg5Y,\"��'T\�0_��а�u�$��]3�%�+�g��9@Q�g���A'1��*�X�Y��4[�>��#ȕ(ޚNb��}譌�[�'2Zk�DzzN��Y��MH��?�8���e����M� ��½��It�-@�h�.\����?�k�N�|��QF�_�,����C� �����fx9s�-U*��h�3 �L��3�,ޱ:�cu9\�D~��	����]�z�b�_܈{�ϴU=R	�-�,�Ɛ�W�
�-���UZ�EɛJ�n���SH���P�{ҩ]]\v�'� ���Gu���? k|�e�}.��ا"!dC�(d���|�V?��`L��4=�S�L��z!�b�<�F���0g��'�a���Z>К�\�i{]/�S@�%�@��D�l�v�ۮ��k2\���ˏ9�IД�\���e�N,�����E�!����wXXi��z�0��NS���w[˩H5�\��P����ɒ�4��Fj���(�)`	�хo���7+^)�j�q!�l��#u���T1	�1�{vL������BH�Ӊe���r^�l�%zw�c�)ʈ8����3Կb�5���`g�����c1�Ghr7(8C^���DCQ���h�&RK�o��\.�M�F*��P����q�� �":ь�:{yE�k�R;w��T�BN���|��o�K����w��*�M9=I��P랤�q�e����8Յ���� �'VT�V��|���m���C�$(5WH��:�+6���5����:����7Cq�p�;%5]��eu������a��v^�k��(k�K���0�.:�%.��{�^^��<�?�;�(��z�2�)E�3ݙ�c�o4�bt�'zlL׆G��ʤd��n�h��}��Z�QOgvuY7]�;0��
I,{�l��w�s�0ǻ��6!FmB`p�����*����v� 2�g�p�τ��v>���^4�K~\6��Mf�����3�Cy88h*BR"ZvjPM��&f�������Z��O|�S��P-c��P�>p���r%k���A���	���Aɇ{S+�5��U��`?�l���WR+;���u�w���C��X3{=��5��p�]�����T����[59��W�Adt4Th˗��S�6�����⽿u6q�r��(��ɒx��zF�>C��͇>�~|��Gva��P���pq�]X��QK�%<oؾ�5�d�&��YG�O�ݐ�줺Ȉ�3!D�;����YU��쪻�qI��r��-_rz���n��H[5�\O
=ձ���R,*Q�cM)��-x�5R3A%��r6V7u�hފ�b�b���� ,Tc%O�3�0���=�x���oԅ�y��@�ؓ�fv���^����V��SI�OzP���aH���k�Ū#�&׻�U7��!�w�2�� Z�MI��T�h힎$����NX�+)�9|5�U�[U':6Pk�Խ�Yu�7�;t%��O�kbx> �)��#�����;���{kY���⁉�o��D�A��,V�*��2�ku��%��]�h��mˬ�)�rC3�鼿K�v��)�>�|��׮�����>K���Lo�<{ȪQ�C���2#4�9�ڣV'�A�����ah���ǀ���^ס޻p�B\��bML���1o��-���a�;�;��֗�Dֺ��N�Rw~-"ߒP��<v����h���8�R�r���E�;�N��>��iZ��T��wN?��w���c.���ٌ2+T�ߓ.���X��:�.���J>�9+q��B�p����"0�F�d2�;s�9S�>��.�h7�?�H�$ͮ�p����g.A�x-�Y$���`u��f�F,��XJBM8;��M�s���ֻcM�)�HY����������.T���{vʻ^^U���1g��"j*h�[��h!��U]���;�����������#�����+_cc�*E=`*��c���'ۥQ�T+v�#ʱ�(�E[���<�����S$�>Ć�ͻ��%��}�j�~��%���Ӛ<؜Z@�X�D�n���1���]��\��,�Xhcq�� ���h)��ai##P���no�S-t��qƭ��rx�*��Jm��=�El̆'��J K�7�^��������l�LD���%�Fh�s����lBǻ�6<���������oB�՜��ϕ�]p��u��Iiw���X���=���+�@� q(8�t��̏����U��ij�yR�����\v"������B�+��٩]�
bO~�]-5�W��K��ڬ;��;u�sr6VVH+D� ���~*�����wH�K;Eٲѝ�9�(}^��g	q�:؄RNzc�6� aN���P��@}��>At��!|��.Z��o�}}���B��S��)�>1�2���	]<�tL���V�n�F�������Sח��(7	1�Q]��<�)T����o!��͢�ػ� �U�k_ϸ��9���1so
�CbB$%-x&sb{*5Wgwi�}�������J���!g��y���ꮞ���֝���<F�|?�ɥ1]��Mu�`C�pxv&�E�]rz��tVfRO ��qgWW���`�]r�HubG� �[t����SI��5^����7��u�e]0߸����X����	������BH�d�A�&�'k:v����6��B�-,��P{�32�.\�03;�fe�s��7��Or��H��ܢΞ�,5~����f��H�.��m|f,3P!$>�el��-����Sd�WN�(^@	������$1/ys��������[l�S
�b�f�}��2Y]B�%R���^Cؤ��:f���LJ
B5�u�t�A��C��Dq8j��N��b3�PR�w(�>��u���ԯ�Q��=KD�����<ۄb���obUu��j�.����´ֵh��kGO���',-��z/xGo�F�q�������b�z�f���L��WF҈>����DHrÌ>�n
�\�"Q7����1��>�7la�����d.�a��^��tIH��x�G��V�����eG�?��e����3S2����Md/	nt�E>��|n���?�4w	3�6��F}ԟ�Z�-G*��R�N�����CX�3u�i�`��d��|2Г53ە����JҍL��QUU�B�����KO�n�X\�v83U����ח��6��;�iiD�B:9��	��U<��p����	oJ`;�u�jQ���[���~�mиw�=��Y��)HgR���ֹ0�j�K
N!d�FM�	��_�K�^ M�D�Hf"舢.u�4X�&{.�ѯ�79�i��掿���rc�K<�Pp�:�|�� �ŝ�@{ߏ��5Y�M�kw�AkJy��<���^�����p����|��[Ӧȵ�[� ��v�?��B���4�h*�j�?�,��9������P���e�%T�{}�����GKf����!�Tm[ՙ��m��r`�U�(���4O�J�Q�ۙ�[�C��P�����b���}w��+��<y8����w�⺫9$Jn�篣(���S|����;9_��s�y
U����:���6 =~��^�޾v�S�=M|	�h��*n)�Z��5v9^�ﺙ�K�C\1�>4mţ� G�o����{�X��S�D���m�7t��U:����Qe�L&�/�*��.��>w.} <آ/��v��W�O|�'1<����G��� �����Ҁ�`����&�;�)����ڋ��������h�R=h����Js��JO ���E��e��3F��?��v3��U�����pC��[�*_��D�O�wۉKh�E���"i�_,YCE-��^az�T�h���Q��eT�"��6^@��sor�c��@��'�1��쏇�W.�(��/j�x�$?��}�V��9X�2&����jv�o1ﺑH$�G�S���^Ȣ:Q])��/�a�|�⑈� _��� E���*�i��<���M�+v$N�{u�<Bt��48I����n�@;@�I  �E9:E+���,�(_,���5�����HO�����ϓ%^bQ�KK��
���CT���C�{u���m/!�^�R�h Eh��\_�?Y�����s�<G~\��2���-�]��z���)@�Aiii��_C����ō������o��>6�<����8�D7��V"d�.��kc�3(���U������z∫h��[��P��P aL�y�� U�o�tU��˖;Lј{��+,�6�p��6�����������򙁯/ٖ߁����8��^u��?�^���[Z��"���m�{�x�$���p�H��b)��Q��A7`OP��e��d���Q�v��o ���[&��A���+�gQ��y�D�G���
|�(�o�K�NļI]C�bgj�4��ֶv%��:p��x����a���ۭ�v���q�:���'��${,4B�.��?T�ڟ���;���ݟ��[|usf�Rl��";?� �p�^h���V���i�`/Y��호��|�S9�(6��ϝ���*��
ȱ)��`���7�y��������l��b��^��ӯ�g�V
��C�yh[T���\Q{|G�]�<����<���.3Yp�$"�G16t6������Qr"��є[-ŏ�'	�i�q�@M�~��-K_v_��E&<]��6���<�@tdDD��fDDtgfn���صޝ򿔚�@�fs��qs{��[j	\,��ߑ�7+�S8{�>|]�9D���
Sg�X$�e�^
C���=��s2���
���N�bI��:�O����W�� � W��7��{Ac��I]vx��4*���'���Ipk�e?e�\P����JL�E��ܟ��65�B��96 @hv�ڵ�ƹ텤�UwY��� H�̬Z��m��'Ђjl��ӫW�b;ө�C��ml;nu9!>{c3��<�N:�rrP��Y�E�.�'w�Z���A� ���H{>�:���ּ�Yڎ��\��T6(�/֓y\:� ��,ߩ�E/��'��nw�?�vtqq����OV���Sc�����j�3��+}��(�A��"��H�R���Ƃ��0�z�X�+ �wp�0=�_���`� ��E�2����}�o�|�!嚹��BE�P˄y;]��N�>��.	R}�zݾjo]2K�����@�0b����"�6[�!��o)�*e�e��Z��mI�aߋ���n��aw=v))����!E@]�s4�z��}1	��ceS�8�K�R콿sL;{�ꍚ��Z;�S��M���۝U>��(N�մ��0D�%|���ahz������Fɇ�\&##өr͓��`~I.�z7tR��{�m�TK��tL��s�/�[PP�b*	Y�9"jv��xP��]��T��L`�T�r�y��9B�*�<R���g��@w^�bB{��SX�|��U%"��:�a��ں��q�5�O(� ��t+��]�wsg�(�7����E�b��'^�1 ���`��0+�+Deq̰`vd�D,?s$%v1`�C]�P3��`���躛+;�
Z��m�]�� ��.]5�X$v3x
�f\)H_�yU�,ɋ��o������2��f���hp,eT�xVb�^>ߡ�����D�7;T���G��s�.�"L�����_�I^"��@w�@���R(���O�c��hm}Ü��2�X������^dԏ�(�Ϊ����D�R��G�n~����YH]���Wd�c�F�!=&���r٨�n���L��$�E:�!_6�'��qOp��ODT���p��u����KLO:_g�"4>}}}���_i��9�`V��? � m��.~�F�P��v���h�?�����!f6ڠ��P=s6�u�eg�H�K���}8`]j�%i����aI�.<��$Յ��Er�&l� ���e���W咥jl��F[5\A�4m6�X\Ϧ��=���S�I����l���<ݲ�*�]����S��dg�P�U@o��F���x�NbF�G;݇�dӝ�l�0�Zlʸ0�XK��T�G����JIF�� �}���n�@����0�0�hɒ�eJ$af�����E�"���;��R��b��a[���,���[F�U ��Ӓ��[N�D�g���w$�&�w����~z��m��0]\��Cx�^���!`��Ȫ�R�Q��P��xC?�I{,�(������%�F�4���"P���Y�(J��������] d�\���mFkk���g�s����e�`<�#C��u���|a�$j`��I�;mU��	���%?��i�qý�B2�������>���{>�j�+;�v6'ͬ�̬¯aj��K�{�C�����G�z��9c�sz��tR$�Ɣ����ܦzVZL��,Ӧ�Z�g���&ɠ��'������N����Nv�#S�.�ZP�����2�������j��Uk�N�P�D�L�BX߱���ή�}�9Z�C|��p�o��T��m���h�2v:#�b�zM:�
��*�kS_nn��ϕ����|��I�?z�^��iw~s܍��]��zz�6F$�^�W���������;�%y��*��U�Jm�V�Ӈ���M�W-���(��/����<?�ǳ�O?��Gw�QM�M�e�OP�F�s�q��%Jҗ���]\0r�;aؓNf|�!�AAA�ۓ�%ƍ���ŝ.Uh(��1`6�@���ٲ�}:�6�1�%����n�F�7���Jɪ<�bM� �������^;͂��m٣�v�`+�I�4��/�}O�6���n��i����%�̴�{[g���j�����w�M�Ug7m����
���Y���7�ܺ7���+�7��7�ݒ��I
�~k���Io9����\����X�)"5`��0���]�]C�7�N�ul�肐ڔ�'&���
	I3a������R ���Ɏx�*��9�W�И����'��/&m�P����:iMp]�����4j�Qt_�Z��9�
��3Ԅ�a��S\&I�o�Sۡ˹А8�Y)y�zh���<��f3�ÇϽ(C�(��e�1a+�o[5/�����1�	JPpa�0�����D�<�9��D�R���1�]�q��A�V���s��,�\�$S�<=noTt-��/��[��3��B��d���s[5�"#�o����)L׽�2D�ա#�|�S
�-�R��#k�(�!�N����gTxyUq��9���;�oO{ҭ��$A���d��0��}vYM#�+�ڽ�{muw��ʭ޾~�켼;6��sH$���y_A����ଜ��w56C�.}j��Z�5ka �.	X�,�a�.P��6��Y;:_���ŭ��-+�J�g���J�ī�f��ҁ�Aے�B�3�vRCKW�
��-���4␰��3tʮє�dJP^}�>n��`����_1}�+��
e�(�M۩l~|����u�5j7�p�,tL�%�9,�	���⽖Z9�_�$%5����ɹg�n�*�g� /���w�JcK������<�����CZ��[��b�>N M��x�nܹ8+���/v��ʫ���F,�^�� ��cϜ��*�A['S��֚v��|�� T���?��9Tf��\ǹ�~F==}���*�.�8@L�ڙ��2�]��˚3%b}տj9Y�_���%��y�hO�4AG��=4��ϭ�,�?������~�5�`��q�F������c�`�}�:��s�{"�k����xl�^z��2��!z��zP�f����Ay�>alY�<ٕ�]7B�r������CϵCP�~Q��Ss"�;& z����O��\K��M�\-nF�v�6��J]έi�A!u�����F�UyYB�1�Y��.�����P8:�`�G�}`�	�f/��_i[t��s�ٴ[>Y���	�� ��uɒ�����rPx�R1dh�h���婏��ξ�4���}%�6�Y��{���gfg�W��~��6M����#/��\l�U
�T��n?�w�ۓ��o����&���t��p3��k�/h�y M���������%�c3g��`jǠ��u��C����-����Bwj8>1��v1Z�^zpX1^1�.�'CPfq&_��=��3�5~��~��b�WJ&��<ֿۓ��Z�4�����n��GA���Ÿc/��\�ը)�N��~�l�3����-J�M#����Sn*���6�o/N�`��2Uy��P�bb(J�zSQ�2&;[N_�{i�}���i�Q�kw��>��==3�O�2U&��>�>��' ���%�[�j;3Zu����wԩ�˯7-�:�a>���%��2�z4؆s���������?s(������H��A����ý26vg-L�_�����������q�5�0,h3�����iY����?�gZ�%_�.����R�[a�&]�@��3�>s�ʤ���ͤ��*�?|#���ڼ�#7�]N:�Xk��11��$}��t+��TZ��g&o�{�e:r]�;a��]���� )�"�v�?��^O�{�x䢯�Wr-ᘤ�S^�M:�l�ӊ{��<?�0xb��f�ǥ}�L��K{�+"��ν�y�m P[��6�h�A}԰�&��0�/y>84�ު�z�j�#����-6�+Wh%[�.��?+�j�z�.^h[��6�'ok���z��-�*��%?C�<���XS�\]_�S����ש�;D��<޸���<���C@Ƈ^ر����>�*�.&[W�{�E�oy��W�vT�_9󸿓hFӈ{+ii�y(�r<$L|�r�(-�������0Z��9>�6���ћ�#��]ö�]"֤�ڂB��}��Mڣ�K[�
�^{��9Co8�2�:k>���r���=��wf��ݫ9�5��}����*�����OB813��b����dʋ�2hƓp�����װ����@���$���@ww��{LD�x�1#��]J"vix37)����s���P�N��03��;&D{>��r��If���`���,��6��󔠹cW�Swݪ�%�����/#��cC�{l#s'�?{ !-.��'��y��g����v��]:vt�*r��d���S�����仉h6�J�Hb��$:et>����ȘH~��x@������u���RbJ:z�kaD�EJ;�n��LU6�}#�[�eͅV߻��#)���MT��%����k�C�q�0[�l�lrgr�X)Rd�����OfnL�C�Ю����'�V�X���Hf~�+5����ݿR�6��plog_����vxp�؉㚩�_f���#UA'�8�+Q+��L�+8����ֻ�͕�|��t��s��j7ۆ�eWKkY�^�Go�%�U�,�Ƨ��E�_QN՜$H:1��_/���'CB�'�8!���b��]����Ȩ�'�/�Gk�$��w_Oo|\�V{�m������Ì�?�f!��U�f�U��R���p0��KZ*��üu��%'n��u@���9UB�2��c�-��A�Ж�]u5�C٣[k+�Q��%��*:S�3^�v��I3ݩ~�?mV*�*��_v��/_���2�^su�������+g�/�
q�b���J��|�j���:l��X��4t�WmJM�K�Q`www.�p2>��0���u���jd�Aى�����Z�ɦz��M��`(��n8T�^����p�XDf�:Y5¹�0�TP$�D�y�{���ܪ�1p�-��,}_�>���L��_���	�
6&���������@T�1ol	
�P(��U��EW�n*;���l��8������5�t�6w4�:T���!���ަ�%~p��Ю�Ҏ�-i\V�e�3�������\O���'�ő�D�Njj��X�� ����\�_=�5aD����#�b�<]t-��?Qi[O@#߭�2.�缮�
�.o���<��SN7a�X���dI��D������B�(X����fՒw"����ɠj�<��;�����ӳ�]���4fz���C��Y��������t9;����W�Ӟ��=�S�h]t�Xo����m���'yJo�v�]�S^x������\j�zp[|Ջ^G�����nv�ޗ�� yN*]�T��<���C���򊉄�}��	���YN`[�}ZU�6�B���QWos7�y�xd�(z�y!��=�o���
n4.�*�I�{�2�g	��}L2�a��jJe�p���y�~2�q���.��q`H���ԝ�C���'�v�f��<i��N��ޮb$����k��w��(k̯�I���#;�C��o��yL%B���oN,)�k�d��k͊�����agƤt�C�}AI���Y0g���������l�Χng����A�T���a��o�M��XS�^���+'1¬��L����y,��}�a�i`����ca͎[�=�t��s6�4�`�6\��R	�6��`��E� �W��^}������z�ݜ��Gl2J��=�J�ʯ��|��)�W��}^�?H�X����M ������r�qs@o�ۍ�Gg�!m�Q6e"�xcU��z�\O׾�u�)뗽���u����f��8*IL*���ۆ,��kDV�}9=7<=ʸ���>��Fte0�`���Ƹ�6=�ホY@��G��'?��ﭼ-�eV���r�a��P6�v�d�;?�?3֔A#�\�gJS����y-0�]�+�C���?y���yI������|Ծ���;a�s�����i��ժW_Reb��s&�{��M�|T����k�vP8�9��]�xR�4N��x���R�'�0��6sa�� �I$3Y��fC��8��4@O�SO����~siD�ˏe��{����/"VYQ�[J�|���:Rk-6~�G+!�I�s���#4�H�R�K4����$���_���|�I�-ł�e@@�t�s5�/x�mQ�y&����#�!+�U��iaw[�N$�Q2w�\�ZV��p�1 �ڦ/?j�p��'X"��N���[����>����{�*��}�xDiRB��PA�D�tw7"-� ��{�Hwwl�κA|y�q�:g�1���ϡc��{͹f\�k��֣DE��f�3�eRp��l��nM�OAzx��P_ʓ�+������|���� �E�f�ա{�&5���Q�5p�dP)���ݽ��R���,�*ׁj(�@�}��c�sq.�zx�>f8��8[�ᢾځ��oV�fR=^�C���4�7��B��?�m��V�7Sor -,�*H��	��{���P+*�Q��Z8�_�E�����>+*���H�	�ߦxJ��O�]Y��7� &���{�D2��N��&��;��ٳ�/�"FC����>Ɵ�N�'�$N]u�xZ~�q[ߖ���(mS�ӕ���F��Lh��٠Uwö~����ڒ���V.���?���̹؟�r�� �N��W(����4w�����A�TE#�}�|����qO���n�k(�濂r����$g�K%�����P�[)n�t��8;��!q�3�&�A�j^3������*��˾�݊-bV�I���d��r�(G�q�X��З*m!��J�P���{vP��-�P]��j�d��dH����I#z�P<��[;��J�ޥ�u��j|�y�+\q�Ml�_o�?>�P-��*�ai�8�����="9?@��$�mI���R4!�b�4���VۇV]��{�O/���:f����)����T�d�8��[����*M��O(7���2m��mt9�h�R�D�� 9q
 |>�xd�C<6!Qv#΃J�|�i#Մ}'��k@ۼ������ǰa�|'�*J��L7F��|k���;Ʌ;^4=�蠖��������I�&�����&'Z��ҥ�|)$�z��U~ h�=ܮ\�8�r~s���5ߖ����W�x+]oA��,��.ETs%(��O�9���H�)�
�-�۹%��1%�rBZch_�{͕8�Yˡ���-��3� ��s���� �mo��._�Ů �� ��݅�R�G�����ғR�(D��(z���>���%Q��X&F�8��#�|�� I�����G�}����U���][��R�i7Y4��?�T�%n�s�z`%��_%I����p��6
jm�/�����
�ՙ�mDH*�2�y{R��QP�`��=��(�9+�1��^d��u\s���/p�׫�0�*n�6������C��g�+���й���@d�a��@���:-�>q�~1>O�n�vm�ɚ`��@�:��Tv��7:Q>��&B�~�����S&Ꮋ�1������OC�xr.diՊ�O ҕ�� l���!.��+�|�8xԸ�zl��3���ťϧ"L 'T����̡21c�� �=��0o����[wvϖ`RW:��� �G���4�Eq������K��˨>�)5�����F�n�ҽR53燖����]^���M�w�#����zH�-O>A��m� z<N�T��4�L|�T�]T�)]R��MC����q^^��~8(+�ֹ����u�D�k.�����l�'��>"��@N�o��"�d�-ǖqlW�2�A���n���h�^�!Ʌ݅X%���{1�R������FO�wv_
��5l���o7�]qZ�	�4�s��`o�TI��U��w�|5�*w^>61����>���	���C��^�9��Jw+����d�t�u�"8ˠ\�`��@Vf�Չ��^�"ǽ��w�`�#FFϝt2���K��|���l�r[�Z8��;��ڮ���s���4�0�١��W� daD�W[jU M������:����NB��Zg����k/������'Gpb]����z1�� �����u���=@k<m��kC�d�A#Yv�κ��O��Vsa^�ɒ�����_E�� �㪖�)
�E�\��R��a/`Im�̛T�e-�X�KUrj�G$жg��M<�4�#���Egz�J�KOLL<���*��d����xĭ�80�u��T	��e=�Y�ό�/�"Lr>��%ut����y���yl�w]�ߔ]�K�Qq"�1ҝx��E�={�{Л$��^e��^'ͦ�T��Y#�/���FW�cG�+��]�zI��2�,�@݀D��Kw�w�w�L��<�ЏWo�&��SY�9�d���R�D��Ǡ��q�:�7�������������B:���`���6��Q�`I_٧�7�ˑ9,#Kj=l,[Lj���E�wP.�g�����`�M�N�!��l�xضg2����@�"�g��A�:�"(%M�M+W(���cM�(x�⹇��ꤔ�ƥd<��e��r{ƺ~������s�
j�nv��	ٽ���sƺEF0w���,�W���*l�ل�/h.�����ʎ6[��gC����@ߑ��6�j�U!�`�����ׁw�
y�g�~���'�B���GOL�1<?!�_BVeu�=4��7���ZDA�yD��Ź^����gӮ �޼�js��s��d�ˑ���:w���|ҭ�r���`v�I9�]8���r�FV��������QL�>�P�G�h��,�c�u��{(6K�{/}���O����>]uZV��^,�UQ�}�����5t�1*�(��5q3_V��D.��;��Y6�4�Ԙ�ta?��Xf�:d�W���>�4�|�~C�Fg�3�4��ڼ=S�Ł�4Vץ�Q��:.���z*����!��~���.����}P��t5k��$�
]��3���8_I*�.��"��ѿl�K/F�>ܾ-��9����JwI������oee���DZo~���92�pKū0��ن�v${qc��[>'��nC�@���ݱ��l{�a�k܄�<d�W�r�=�wz�G��8�x9	#�����G�^+)E�2����dE�zd��[	�
4'���W��+�(2�^��>��t���M	�T��n�4:�Դ�ļ�#��O���	w6N�չ��_i��ƋNSo�#z��e:^�g��-ah�_G�=�-wZ�\r���:��S�]!ϊb</r+��Iѱ)��K��h�/�姊w��_��"aru+��Bկ���9�\�ey>3����%��re�.A�蕷-Ж����U��u����0�K��B����W=l/&��yv�u��N��}&�p�٠aw�kB��h:B
�%��Hz�og0�mm+*�>�:jE[��L�&F��Q3<X@��M�Sg�U�n��t�p%:��r��i=ZV��?�=�C���E{�Ɖ:��xQލ[T����5� -�u�'��4��!T
��\�����M8�w��?�1y6���Xn�_0#ͳ�k?P���]��|��DD1���t|�5w���"��_n}r^�G����F���B=��Z�t�4�d�g<�t1�זw`)J��N���MT�ろ����$�Z�u('��A+*���3�~J�:��G��{����*F���0��'>�{�������F��l�ѥ����֫]>D\ }�D���2�F0R��`��E$��̱���ɸ\[b7m����8��.�r�m���\Nt�o�we���P�ؽ1��;��1/糩��r�bw=��ֆ_R�/�o/�*�Ď_��f���=##Y���#�Uf8�5t�:�F�U��]F���˩K4�u�6��Ҁ�j����ȿm5��RC��e)��t�+���	2�!�R��"��s���B��$n#���b:��?�]�}dr~�	�k�p�Z��")�&= �}��cATis�\�6N�p�M�#�Q��-1��1��T��c��D�S9 �~��Z���[n����-�D�t�.�rT�\.��8W�3�?�x���GZOP���=�hn�3�kW&N�Wx�mf��|��̰L��s��,,�V^/�=��%'t��K��`��!C;k��1��T�ݳx�bޮĐ������g���������I����N����Җ��B-���-٬5a7��?WϿ������[$�H��y+=��>4UL*3�[�V��Ͼ����f\+���WX��</(�Xb���	>45R.�-'-/��7�&x�Ԡ�x_��#*/e`�1�\o`���]ά�_K��uqxQZe�&�������S$�f:�֊v{/���#��ʗ�A>�)�"���jŋ��k�s!�B?oYa40z�J�3K���bQ
G �Z�db�c����D�7�Z�}K�X!�	����WAi�f����~����1u�A��t�lJwJ���[�^��z!�z2��F��;q��J}ͦ�-�JV&�����_l�|̀�^��x�P�:�/i�U��Z!�j2��O7?�*$	�-��d��/�抓8�:ԋ	-*������æ���B{=<�Z��rWM�}Y��q�[
& ca�����u��~�c\+Lf�8vb��~_�f����nW�{� xG4%�ٜT`e��/�����,(�7�����@�z8�����yt�r~봹C���o5c
�͝TvmiNM�?�@4����-}{�U+�~7n��%+W�`F���i
G�\h� ���_��B����䟥���=���F}Ez�H﮾���]��d�j�d:���1Y�I���h����ʬ��+���/�\�l5��؝�k�o��knk�Y�O��&���C����{mk����x���r�hn��vQ��Q��������Ğ�A͆����!J�:��%=%�_ȌjZ�%Z�>��hQ��u�����Z�x��:P�����T������J���6���I4�Y�ae��7��7���"�����ԭ�5�:
4y��hWf*���z/�����s.P�˅u�$�DK}����%2Z%�aB���8H�\���M��EɽP�e�4�Ӝ.����[�;�\������]��6$g���X�)�U�S����?J}�9���[����G��֜�h���9]+�ټf�f+��=R��~����[��.J��t�(�΂�]����vL3֛x7K�td��ʨV�Hs����ʧ-��\�<1�v�߲�|�ꂯx�g���*�|�IG��J�;^� ��uP#�K�]�쮔6�;W�F�u�uIE/tz���~�hjhm�u;,�xI*�n���L�|Ht3MC��'ԝ�bb]���)Y'��ģ��Y?��;t�R�I���]�^�
�{�G+ŧum�޿`k2���U��6�_Oߙ�K�I�c���2v��EaJ,���|�8�6�|�+]��+�<zQ�����'"	4/�M�C3+S�O�+�d>Wv��@'q)F��p�l�$jQ|��%��x���;�n�Y��VϨT[��KO�>�+�\1�5co�����>�Z�A;-D]���\�9�&)��5�lP�5̼0���6�&`L~6b���M�Y�ڷ��o�Ǭ��*�����a �ڥ/��F�?.�sm
/
�"PK��ӐeC�N����P�XD>J)�� �HVv(�9x�k��B���[�w�=��ȏ�Z���B5�W^dF��8�����S���~[RekS�yЭ�tL"�-zX{�4{;��,����t�[�pX���Ո�1G�h�:{�o���<I��2��{+z��9J�G�ǼZ>���M�jw�
���O��	�d�ɴر��B%�.�v��:u�\���4��m���w��G���Y�:�?n���_f^�7�MGU����W(�댻�����^1���J�������~LN{:��E���g�� Pnt/ⳇ�`�u�>���[�e��^���ֽ{�V�����������F�QYHȆ����K�T��yC�Q�[hQ'�)�{��)�x�h���{S��T@�R�q�[yB�J�����J��D��4�W/N���k�Vӳ>꾚�)S������:����PKTJ�����Gۡ�Q�n*�;$�+��Oqt�W���:���V��+�j�9n�OLm�������!b���Z+=@�Sl���D �ќ�_O�r�`�b�����3�{l
L���v��E�j����Kȕi����I+��Ϟ��v5���wI\֚��Q�+ӽ`���6�zG���F�㳫����H�3ϋ��G�h�=��G޽�c�7�E�P*<H�A���6�/�;����՗ȝ9���fg����
Pg���&�65���6�t9��y��W}~�?�� ~�{��`�4?�y_
E���4J������Џ�/���Pgs�-��O϶�d��E�s�s,+�u�Ie�����~cR�N�1��!yx�1�a>�?v��>�CR��D_�=!xQfd�oG�2���2���Z�A�������c�D�櫚�]Wq�	��xSI�k.�c��)����b6�v%?#
f�7�#�2e�k`n�/�5��2�_KG��";P�)�עB<X)r5�,��9ʘ�_�,^�Ę�#Mi�G�r�����:���}E?�1��G��%:�c]Yo]��5S�89Mb@ܬ�?S.���_d�^�����b���P���9/����uТyJ��0�8�h0f���F@����n+,�NQ��cT����?	_l1~4��Aρ&۞��gI��p��c�16wi���n���\��#���5VX��9{�d����-�P�,�]]^�$�T�T�`z��Ov�CD ��3�՜t�\����] ����5�E�t��ѿ�<�S��*��ʿ�a��A��y�'���5k(5הvuTй]$J�V$�j�{Ǽ�n�hnHԘ{�p�]S�)f���elq���_f��w�hk9���1��6Q�����gM�E�8�m���an����b����w�Jnהܖl=�����Dk.d6�;7�M��V��-c"�2ܺ4�v>=C��m���B/�6������u��mّ���s��LS�T��㱊�p����G!��B�����E�HeI�'.s!Y��߹��&?	�愈�+w��%_o��ů��b�/�Ɂ��GY����5f2o���L�9�M�a7��,��w�F�W�ȏ����:�ws��>g���Oyʢ⳼�&�o�����VU��ֲy6�s�_']r�[L��.l&ˌN��]�y�͡��p��	в2\�e�������O^�܅d[n���.��XI�J�>�noP�W:�F���8v�0eT8Z�L��&�|��f��Q�w}���?�\�Յ"#������:���<㿘���5`�_�V$Q��a}��N~�x�u���%0!�5��ȳ�;n^�d��GH.��?R�&�w'�1��^��U;�يDWP�&3Q�~'����,��O�I�R����J�ճϥ����>�ndxu;26e��)]l'3�q�������*��a ����X�s�\���l�U����i��\�>y}�Q�u�[<}�)[r!Z���2�gv���Ꮎ{�CKp̩a����g���-��Z�X/�Q��ǵ�_�&n��6.8d=)g�p��/F���9�8��b������|��,!|M���)hY�����x��<�u�	��z���gA�X��R|/�Bwd/�$׮p(b��{��㋥N��lY<��ao��N��{-���;��v��q�D��x�f��"{x��-���qՃOvz殺��p�1PD�}��g��ʣ�lo\�����]����8��TD����]��'�J_���H��H��Ϧ�Zs�����-�+XF�+C�e��{��̥<6��=���o/�����%��t �����	�#���OU~���@EA�*3�J�ǃ(&���rK=I�K�'msGGW��|����O��p�K�<�n �^&q��c.�8DN��|�r�o����R��pq��x�>:p��N|��H��t\�>�����i#�?��x�"��n ��!J:���˺^�N?�P�2:������1L]�(�q[��Ӗ�o�\���ϡ?d��e:t�%"��2#�f�U�|_7�?Yu�5r�c�����H��9vKr���^��AYxV�0]@��NM-w�^��nUݴ�f��YW��'���q�����+st��p�����{4sn�к�&A]q�J�<�R�B���ZC5���^����M�;Iנ�Y��Ĳ�O��7�5B���r̠���b����� � ���fg�J5q���Q���Ox�,h�� ��jq�%��;Ʀ�$^�8�1\�C�h<����_���f�bJ�6)������g�X[M�l|:t^��v~��w��%'ǹ�2:<�N�q��֯�&_�}Ǹ�_��b/�\��җE_+��6m���?Q�_�[��2P3{�J#<�o��m���5���W3��I^�#}��p�i&K�U�㏶�����s�$����5CG���*�l��r�a;��*�� Ԑ�:�)w��S�&:٠��!�g��lH�^w��m�rF�v�Pٟ���!}�H��*�S�8F�=����˿�9�Y&�:"�^�����{��p��p͵��:�I����7X]?�
G�Yu�Z��$ߔm&�Q��A*q��A�t��4�g�K�k�ی�S��-d0(j�+����//�T��J�F�nR h�(����&�@ި��Mb>#T{o�2K��6�1~�w22s��K���2 ���_��})p��ŭ+��&{�ĪݍWm�Z�,'�a*FC��F�����蛕m��t?���F���v���x������-wǅ]W��hu�u?��.�����G.c>��mC�`��|����D�bǌ��ZZ���<q�|���<�B����O��WH�d��Y�HA��2e풊0Q�j튷w4e�l@��շ�#�+u�k�z[����tkSP�	4g0v�o3ߩ8����M�=�Op�~D�
�ct�)��1�ISOG�8l�ՂS��i5A"_\���@�Jo�2��( u��}�~P���M���g"'���&���OƢ!U)�ChWԾ�}��owq�ߏ����?$
B����A[�!_�؎:�c�J�����$u��������y
'q\4lw&z��bR}/^��E���2�馅�Э����O{!l�<c�����Rs����1�����f���9#GU�)������{c#|�g�"w: �|���m������zL[G�KI<��:F)�3���?2Tc�T��Y�f^��x\��$|k��Ỗ�>I �p2
|�v��	cg�cy�sP��;q�;��~S�o,E����a��NN>DL�"t��W�x��*܈�q�~t|�m�6�����.�A\6�M�6���.��ŇD���������%;���YHn\��Ҁ�,ϑݝ!�� �Pi�$���ѽa#�zL��YvÇk���-���0���~A��>i�-S�V���jP��ȓG�c$a#[���1)�5�گ�?i���.-e�~;n[1?M�����ƌ�0�Å��{�wFg����H�x� ]�X�>f&TW�UjSm`ypT�?zͲ�oӶ�J�7��K��Cou������y��3wT���'�&G��Vq���𴟮.2��V��x�����$���W3�w�4�@L<W�b;��~�mD���DJ����]!I����`��|�M�F}�����,�����ʠŢ�[�Ю,�̀'J<A�|��%
��I��'hǉ���W��D:|`ǵ�+v���|�_��/*N��5�'�	�?|�K-��?���{{h ���D4y��������9�y�Q�걀��=�X�M.'G��j���#��4K���|L����p�rxr����145-� ��V�;��JV7���%�|�"&~zե��d���]���>��?h5��A����J����Q_�нD�*��.���^�H�B����W�ߩ[�M����\8y�l��uT�5��6�H�I،���0M�ci�7|�x\u�YO�N,&mR�0��m��U~��
��E�)S��zU'�����E.><�y����>���x.��w0X\�f��:`\lY㇩o�흓��h��O�	�բ�7��G�����qc�E���@aܯ1��!ݼ��������ezh��-#J~��l��mRKL*>��Z�ڦ�4c6�%�<�8s�H��*
%j9�''��*��(�Wsbb�X9|P�i�ҚX��wb+N�z|2��ʕj�ڤI:v2��73�0]����q�s!�Wz�yU�8�K"�S��uVz���|�c�E�R�
j�4y\|�cG�[յ���P�����BGR�p��� 3fp�d�t&u��,�;c�@[J\��,<q��ۍx��]�|�]�{�λM�����
 r+7fR=���
��I��������v�'�}�p��=����)�I��}�S�����&�D-UM�ӪvڲZdR��Ω��H׻��u�A����'�"����̑��t+��e����P�lΩw@����v/�.�����ֿq	JV})�
�4�r�
ް���LR.Y/T���M�-I[{�e̺W�my뭞1��)_�*�>����a�����\��4ڲ��G�llq�|R>���<��O ��M��d%-`���k�o���ިD�/��������E��p��s� $S��T{���+��!e��,�콡��oD�|������Gl���+v�}�y���)yw|�y�W���r
�zK6��;P��7�j��3�(zhD�E���r,���y���qc�i�*&f�!�C�r�p���.�?k�U��;کQ �����pp� �xo�;�=ض0�]�w����9�� @���;Ӎ��7�M�T���Y�n��r#{���˥���N�<���:利��Mۑ�̱�P���e��oR<#�տ���;ڶn�䯷�S�r�h=G��7�L�k҅��ި!3���	T�c%O%.U<MXIO�h�7&d��x��h����6�*es�%&q`��H�<:���!�f3A;ejF�^՟�<����a��Qg%��T�kUȬ.d�mS���d��l .ž��!�+ĵ@�B��҇$����o޳�2��J���0DF��R=�a^z��a���v��.#��������6���q�{FK}�����aLiNM�p���Y���n���+�gAA�����B�ܞվC�ո�m���p�⺫�G3���2��?g�<V�ғR���[��!;��xE��q�T�Kt�ם���7ji˪����3�Ucm�����B_��:g\=�S�������)�z8�i�I�;O�v:��˂lc�צ~"%`X1Z[���>j�[�a�X���]��|c�{�ޯy�iO��������0U����n����Ķ�	��v��Z�s�_���jx�]l?��KB�m^q�7u�p��Q��L�VZ'HW��}�0� >ݿƉP�����r�l��2�2`��O��g[6,�������i�Z�~�s��-�ga�\���x0y�Cts��/	�/1�]o��)x�ϝ'?i��` �������mn�	M>=_�3e�v����)���jۧU[H�����������6��w�U��-^&V��B��Q�m���q��S�7�x��^��;��Zx{�� �h�y\���čGR�.�%U��X^<��k�^��wX��t�M��ȳ�t�a讅��<���b7\׈�]�r�t-wo*���J�nV�Ǧ����%�V"*�Us⧣iX:rF��1T��ָ����rZq�Wg�Б  ��2{���7)��:��hat��zݣf�d���{�~:�8CJ6��1�>�=�����-� :	���g���AB�q��K�Ҵ0`�8[�W��IDJ��d=��a������	��\��r�D���J.���v���i�������3ri����g$C�R]>��ε�K?L��_B��,���.�#�aa�6U[Q"Zڣ�B����@⵵���sL1"��v�U������
u�L�������~0~OJj�e3'�j#\���7��!�'C�u��t�H���{?��τ�-�_2a��H�|��j���t����+SAm���g�������L��B�?��
�]'���HsK������z�۸ꆆt���{�C�C΃���ĄUYY)�qI:=���Ͳ���/�)�O2��
�_��+���?�
/��������쬠������+�z$�R\J������~�f�J&N�&��?��L����ה������<񎋋{����ϟ?�K�Q������o��_��צMFJ��Ƿ��54�588���������������I���ӭ���Y����< D�P_600P@Mmr�hݵT���W1Zfcaَ�Zw��۳}_fI�T�����t���W
�	��%%젢�gdЉ��A/���q��_d������d�s��`//���Fa/8xy_b��+!�韮�����CU�1M��6��~Pp����V,��蘒���ؙ�h�qy>GI.�oMk5�H����*�������tu��u%�u���3ps�|�z������y���̧��J�iii=�)��%��]�U�m1}����11$,,,o��dee������ζ�x;�'&T�ܽ+hbb���n��۴+����67���h����8�2�����BBB��RR�_�^�AG����#�����QZ/'��䥥��������5���NKK�i4g���srr����G�к,�UޠaOO����20b�Ѐ,���Ǡ)�Hll,����l�	��EES�kkt\�ƣe���߆��RRR���yx�PQQ��FJ�v!�Z[��)ıa���v��RC��㨵�,�Y¬�#@kA---Mư�'�����yxx�vV���K���=Ʉ�cXJZ��ׯ_�����{�!/���!;v��=���S��i�t�I�lXX =��Z�ÝU��	ٙY��4}�.����ڭ���k�<���1|1�;�?RR�{���\Y���n+���65�:<<\}u���	Z��Ey�O@�v������2k�N'L�90���ۻ�ׯ{ E�������_}}��������A���(�2���u_�nD�VP-�Uxll�#���BV�?*ŕh�v1��@�pNo H��Ϸ�l}oӎ��e��T���HK�#p�]3a��#yX9���W��QIe��\]]s��J�42��ۣ��e�@��:�@����^�@=���>h����N��U��!!�
ڐ��!��!�l���E�,����o���	�?�3����T�56����{HB�����n��iim_Y1���OD��{�g�HYEZ_Ldfa���Y.�/++��ۘ6;@�Q���+�3V�oml�C!~ [r�B����|H��A��H�.��2������ /C!��5,,,0�"�󑭥��@� �)-�FK�ή����:�u�+,d����}������������Tj�d��JK9��G����n߆F��j	.��P'�s�v>X|HD$a��Y%0;?�8�^�OL�XZ^&h"�q,��^�t�y�r��kbb�|qv+
�Ȗ��l���`���>��� <6�qŕ�s��ǿ\��gDD �PAA���E>���x���E��$vƪ�틽 '��ň����q����!111��<
`��h@8 �)q��w�����yX%(�����S9`>DT֫C8DDDf3�~��%�\�_��ZY�h���x���V1].�#��nկ���l��������5Q���7"�4շ�zE:�n5ut�������B*W��N����--��L��6Pd����L��FA�$ �
�.�Ä\�t�����֬�zto�ژSF��Y��cqY�|�M�� ���nܸ1o��=3����A�PL���c\�3x��|G�or�3g��\Xht4���WM�u�!��~��^A8�l��
�t��ƈEǭѿ\b��Sd4���z �08���r���Bө���˘t�4��y󦠨��:|�nZY���-&�Z�@gg=���Elq G�4
�Aap)(��:R+�d>�<���Xe[i���&�Tl�}gu�=�� 1�nSMT1^����Q�����ά���~�Fo�Ӊ���X-�yT�[�����Mf9�uk�T�ah�AA!I(W
t��\�~����2�ؖ�!0�Fo�,�W%�+��lE&��B>��;;֙$�_j��Z4s���JN���/r�&M���Q2�d98<��"vK���5]�8%���h�����b�ń  )�UN:�";�����"R��$�����B�Ķ�l��o��l�5�v�OH]S�|Q�o�xB�ݸd�kJz��=ZEpc�j�0�����?���g����@$vhHRR�s�~dB��挗�倨^?���p���\��j;��i	{�Hv3Rt"Nl0��6*oX#�W������f��xnf	� �")��Ҕ;U�����%.e�F�x�J��,�rR(��C �@����{P�82B����$�AzȐ?|�TT�P�E��G <�!#$d7��s�9��.g��4��c�� X�sA���6�92B�˽)��
�"��|��?AWf��}�J3�1;�cd�ƀ�oCO�ۮ����K^W�
�/�W�@b7����#V�ǉ�$#�}��l�+@����S+P"8�l|�\	� 33�⇻�YYY�Q�=�bttcQ����7zT�i�v��κo���ϔ�$Ν1ӗ]L����l�<���jH�m��s���Ў$IDLA�|SSS	�����@ ��J.b�t>Z���'����@�b>�q��l!�.D�i����]�S�B$���D������*do��������{�g���K�߉m졋E" ��^�����.�a��}�X!-PMVN��H� Y(x�?��x�q�-�l�0qJw��%٦�rA\�_�Ft.<7�o�䪀J*Z����nj�@�ؔzG4hB�Q��@��ç}���x�߶��C��+�V� ��I�����x�?%�}J�۹.�'��^6�' *�*�e)���h	/@<W:��A���I��K�Ni
�r�B�d�Z����f����B��t��E+q�����%�u��*ޱ��������zw,�3Wn�ȇB�-&E�ƵH�]�y���bD��:�GXX�%4� ��W��@�DbC ��0�=�N�~/  @DJ��?#�����{O�qŏ���D=}}pT�{��H]2@k/��'�#�A[�5P������7��A`6o��O̿��?i:���RYB��oee5b7A29��c%�@H��\ۨ�;���.�
ظ�Ȧ �qK�����Gj\�Z���!Q�c�q��|G����eJO��>%�������r�U�Oۉ�7�@�%"5��^넧�<�Ӕ�?p����Y�BSj3q�/!z��,��722 f�>�8�5`w�]�=^>�9+oee"ƐI9j/�d�q�4�f}�*تjץ�,���"�DW�|R��J��������7��{g��7�R;4�UQ�O�+ǋI�
Λk��Jh��f���%�\�Դ�I��O����Q("�'�Rח�%!�S}����\��{҉�W�.W�~;*1�ˉ�b�s%��d=*>>�ǔa|.U�h_�?:�755���5Ά����>2�?vV,�zo7tT~�}�엪!��V�1O��~^���.�Ls0O+�|VԌP��&usz� 5-m �."�����u q�$@���A����4L. p߽�dɞc�{��#�:!�	ӌ1������OT=��?$��`�?"ff��}z�u��Ua�e�PJޫ��f�+/Z �F�Y�
� �zB*����X�u��펂*<�����$�������ԏ�bN���;b�5<����g�RXs�~�-!e��(����'''��2�UX��&6�AL'g"4r����>c� �kl,�:���4��A���^E[KG�c��X����P���R��~����K�+8v2���kn!i��Y���2�?n3�q�{q�{q�g��{�IQ���d;���8�*_��`���TV�iR�P��(r�Yx�"��7�Hʨ$��Ր�����:*a�y�{wFx�������v���^y��f����< �H����7�*출��Q������ޘ>_�t) �Hӵ��NN��й�t����0������H/_�g��&rvP'&�;Y�`��&l����Xd��8�����`�` ������d�+IIY��&`�SҨ�n�&���r��IS���k�V�1KG��hV�l�+�9��M���,t�q�����:��8���Ef��������ꪓ���D"�30���GԛSCF������!:\���'��9}Osb�\�����@�ܗ9��_�sO�{1@6��$�p.���=?%�Ӻ�[�RR���+a�0v�5\?��ݟ.Χǻ���]��־����A6��@�Q	Z��FЖP}������Jx�<ռ��\P�������c�m���`�.��������+ww�m�ݶ�v�[0R�M7�=�|����11.�pZ��4��q�&<���p&H^��������l�C���1D�8������o����AÁ����j������QRR�MR5���9d2h'~{OKJ����ȷ��۷�Н V�Ag�FC�6f��l�_(�d���u�=w�0��d��h��f��o�'��߂m�b8��v%��bc;�?�������l��縒�o\���xy�_��ۃ�t��������&g�//.�1��<L������;-\�2h�~C�P!o��in_�=L^R�д�t
���k��C��P-��S��Kq5Ȑ�	WTVg��d~�ǠR�d�����؆|q:;��:є���}�`�5�)��k��#~4�>}����퍍���l�QX��p�I�ËA
ak]��ޯw	�nvo��ת�Df�E}ct�l���9R�sZ��XvKl�2u����Mp��I��xZ2�jWP6(�m1�n��t�rw����h/i��7�)�������o�6yBOS7�+�,������TT�!�˪��!L�U�lnm�T��T�d��������׊�HI%H�,���<��( p�;nǯ���8�J�=9�^�=�'=*`�a����Vb�Je��ὸ�#>�A!�܁qh؀-1 �����f,H��h<=<N�DNTA����HquRJ����;��v㛱Ľ��w8�Z�eV�!!ɀ��n�� bCU7i���q����hI��Օ~�W��=t OQ�W�	�V�����cqQ�3��~ Yє&��e8υ� ���:zqee$,(h���������xu�������&�.Q�_�vy�� gV��t՝�0�����ifE�0@�_�����;�L�W��<?i�>�Lp�bu$I�ˢ�9����;��o����́(t�B��`jT@�Ò�0��ls��ՁSY��"� �f�u:�V�
�W��w�|	�������C�t������恶�Ʒ}	WWW�6�-L��
�S�Ӈ v�m|�_�,^s�$�X���xy�!,������PP�4��hֵIsS�oHʣ�|�Y���-(¸L*�z��M�Rʆcvy���p�䒯�r �����Nz�{�n�D'�f�6Yi��i��R��[dÙ-��gp��>�/\���1��;��c�1\��y,jb�>l�F�y��nk��5i�g�v��j��f�u����N�P��Y~��U�Г��N�<̉ezg����Ymllܬ�F�K�1����Pu�Y�u�ǂ��y]�r���&(�������_� ͏����O��I7K�<���G��N��H	�$,8R4���h�ٴw%}|�y��3��b������q��[I�2��P��4Y*!D��k�2kc�ne�HDbH��%c+ً��3�g�>_���3���׽1�<�sy<�s^�3�w~D�4��h�ĭz}M�x�2�����4�8f���w���8��3a���m�H�F��t�_����xtz(JK�͍H�P��e�ίc�`�?�w �,��'�̘T�\I+�Ǳ�w�Z�N���>��m�R�`^�4k�hR�Vi�R4��"�4�6�[�B�RHܞDD�=�kRXmS�Y�������8����d5�/�u�%�Ƕ}7�_�\�$��>�ӽ8�|e4�\S#j�R�A��)�� ��6]s1Zk�֪��^y����&&eQ�\<O�H{��F�R_ig��Nt���Q�w�H�-@^*��OZjϐG13U��˔���4"_"����τ�M�G�s9�J��R���:s���M�D��r����=87��\���g��������pj���r8]�5�=��=�3g���IV*�F筥T�\m�SD ̮A�����T<���\�[�=�*
~���1�V}��D%Y��g�
獩(��lCb��H�~��2S�H��Щ�����]�����)
Y�Vtз��e~���B�$� +�7��w�r�[�|���?�̷�	�.��F�2� �3+Ay&&&��q�*W�F"�uv��ފ�e�D_H�,IE��^�����\���'�\��k�O���N}`omkK�Gz���a���9�X��ˆes�ː];k�{Y�0�w�'�ϸ�~��*�L�nQSW�^u�lŀ�;�+�����%���>�8����y�E<���O���=�Z�m��NM�T0jeśM��4�*���a����H���x'�>��f��BU��B�1��4W�����o/oc��g��
]F�Y��4^�J�o�l�������g'7z�TKSp����O�\cD�mj+}�'����)c��q�J;���CƆ�0h�c��!����L$R�.R@�|}i<7�_^�C�N�M�H���n{WL/��@�d���s��f[��FN�CG6عkW���kFJ�K�l.`���_}f���~�W���ȼ��0��uH�/�qp�$SO׷��)�}(�w���z�
?�}��#M�fb��<�g��`�2jaϚ�}2DY�d��1I����s�o�&�K=�T�7&���`]�<��S����� �.��@�z(���U�<4���F�71C��鈴O��� i�?�������o�6��'���<��s a�6�k���A�e��D9C��{6�T�c�#���Z#:�`�onv��SO
������L�|	�y���(^a��v����1��������(
U��
���*QΫ�5�Y�Dk��F1���<����;���5<;�F�7k�R�eJ~��* vuuU���=��i��i�������UK��J1v2���cTMM����ЇE#�)��*���%�� �ԩ/�L�˛
P	��t����6a���p;7O��533�rqz���~�f��k2�|#�J����ޞ������5�pQ0�"��{�9�G>N��l@��1��V��??�J�;�Nմ��">��׶�$�;�{6�o���kvo��G	E}k7 �@ΰn��hr:�.y����vi�P99��Q���-rqȞ�8���|�����o̽B ����:�rKF�����>�&��s�A�7�.!n|��N�Q\g3+]� )A���� lP3k� Y��$��Ԣ�.ʂօ��lq|(�`�4ȸ�J��p��:ُ!۩�Nmmm�>��_�e�n��P�~l���g#(Q�O�>�k
��eo!T��*��z���(��G/^�S��\��i�q�*��<e�R56�d\�o}E�6QSS�kM#sn��|��5�t�$V3I��<�%�Gzz�
���w��V&������ˁ���G���I����F���Ȝ�c�N}D�>�  Ѥ0�P�!+j��5ccљ�殦�Ǚh�6��b)����0'��'�so�
����/�]Ϟ=+����և�!��%j���F1�e�;��!Z8߲��6E�C1�m��C� �����̑��h�r�#_\��xV]�*��jm���E�j���S���u��Y�H�W�5�秉������X]0a�P����8<4T\��7u�f*۶��Q�l��՚�A�"G=����Y�������(�I����OB2�q|�k�7m��45�=#Z����ː�x ��vv;K���_% j\�P'=��tܸ�:=*�<^�dّyc쌼}a�X��טV�-�l;�rY��]����s�t��'�O��ݼ�m�j�d�왟�fU��A+v˵ �h���O���b�a?~��I[����.�x��D��⳶�������ަz�.4|��0�B�|���v
��0,���X#����&���f���p�ib1��B=`V�P�_-)*�?�>�+��2������a�w8��	�g}hf��۫��m��O�2I���sJ�����QBZ�M?��h/���rJ~�E[�κ�4��������'�m>�^v}�kԛ^^u��隚:�yz�H�IeK,����ok�Q��`Ȣ���Z9��_���>�H� :�M-�B�WV������W�DЮ�8�Kt�X��G��/��5�>h�Ħ��$�oBK���(���N�|������BX���DWwa��tB{�e�CC����Os�^�O�� ($��'�!��o��O�U�����{Ё`蟷�%(e�����r�6���S��{��%�3#����5a��ZJ���v�!f���1T�PU�U�u]�Əq��F�(1���x���.^vm�qvaA( 8�7��OMW2�酟��0���3�9VWW�ἜsW�z��{�Jۻ�����Y� fEc�c��j�ܫ",$��-\��FK�tuq( \
t���A�%s��/<�rT�<�����z@�j���V�lcmpo�O�>>�7�|�|Ｌ���v��ɽO�r�榦k|�����:9�uwq�y�}����/PTB}���^ qOV`ۖ� ���	�����퍌G&3Fo{z T��X_����漕U��s�a2gNu��>��l:�P������<h�uC�Omv��m�ܜ�X���ma���1��y��/jX���R0_qL�(�t
�!��ý��au���X�1.�:s����vq�����h#n�˔��bc8Z~T�j�+�x��-���y�`�	% <�I|�O=G�1���	���2�#5�t�f�m�3��W�@IG�d�+��~�W��"�<�Z�e/K��S�|��. ����*,.��D����K�姌��)MrB̇��d�q`��ƴ<;e��㳓��;�*S/EY���2gJ'T���,,gȢ���S� ]H������#��{6M��1:6VHaKjW��;(m��JQ�����7�� ��@���被n�ɳD�&�H~^����u�p��e-["����|P�S��Ah��t��Y�q�B��
\��Ŭ>���,w�������<]?�/	���8fD�Ѿ|�!�k�����w���O����O~�����hoWur�O�$�o5'������#˫KKK��C��>*J�G����<E��h���@W��/��h#��^:�<�9y��{?��^ڸ��R	B�s(��L8�e����x��~q����\74\���6��b����yR��"19��ܵ-�N0Ѫ;n�z�m���*Y�.2��������S���|1��%�����	";�y���y[�J_����{�,N �~�.���3?&�����ud�x��s4ٰ � nkg�D��o4�ܠ�xf�4�W �]�i�o �t�Y��`(��`o]�ZT4�vW�^;�$��:tC%��V��EE��([ܯB6�#̔+D��,*����j#_�f*�^����_cS��S�;"��[�@%��_��ŸFU��6���3�$$`������H�v�f��5pc�����g��
E�h+O<����Pm�4�H�7F[�`ᴐ' g����Ϧ��+J��İ�R��T�:��~ƅC�`z�U���9��|� �C���g?�"˵u�z]ʁ��H@��)a3k�� 9y��g	�\��uc���H��W-䷉��'h���y1�DU,��a�?��m?5<23'g~V���]gOլ\����Q,y����|��V��Ͽb<����Ν;� n�.r��Ç{l���ss.��	)��;�O%݂�=nR�N+7��%�����@Z��$���Lz%�򎓝k���c��S�~d��&�PX���]��fy��#��h��;�����O2<�+rL��j�=����kܶG9ܵ�Ԍ4,�O��Rn4#*�~�^���
���D�ieS�����܅`�n��5���Yߛ�7�7Ҕ��;��^�����_�d��O�<R�?�R	�P�}c�&ƅP=H:�A:P4R��v���т��J�1&��]�%M��jb"��E�K#\��c<>/�v	C����k&���BC��?-�,g���rbGm���c�w���v\\���=��v�<#C$��-��U��y<�;��ˊ�����m�>77��qc��߷s5*x���
aF��,Ot�X�:1�x�:R刬��
ޭ����_dѪ����q�e����׎#�ra��eD��U1���qy�l*E����Xk��L�ɫ׮���[�x<��Q��l��֯UA�I6�ϛ��ǘ���w��#���,��㾇�i���
"�������%�"�Ǹc'l��JI��2��n��q�BU�V�Y%�E�7]d޸ߙ�����Y�N�b�	�/_��d:PDH��u���e�����@���w~���� ^�G�l���E���ۜcn�P ߄~h��2�
g���NX��H�%���M��rU��s,-�T&�"�C&�?�lQ�lN������_���m�!EX��Y��rb��rK�E��k�V�����=J��)n��e�1Kii��89�B\͛��&�������o�v!��sc�J�5���M�\�ĭ�ׇ�^5,<������DWi���S5\�X��w���.�}I͆��111nn_�2`�~�}O�MI-<!+3�1��鴐� �O�2j��%-�f]� �ʩ�f��D�Dʛ7W�/�m����
�V���|�*��`��<k��ړ�и	sp�xG�-�x�%�5�V���WG#��J�����0
��K>��7��i�ܘ{/"����ҁã-){&�ʖ3`_bCC�:1%%E�dq�3Xݖ�y���P�׌���F���m�����k��'����=<�7��a|E^SJ��3�I���2����~�WKu��ڬ��wbI�B��vz��+���`%�`~����d�]��8ت.ޡ���TpL�uI�v�5,Z3<T5���{`P�!s��JS��o2E�{f����?�������K�z��4����k�N�e��",�%��~��2�`��7���V$1*�A�������_��Nbb���ai�{d,ha��p�G� �q���kVa�3��%�a�Ex�P��|MQ�������S:P o�I7,/�+i��&K�Ƒ5�f���_�� �m&md�Y��W�N �J��X�N��l�v�����@�,p�$�VVV׮]{A��ຉ�Փk��*�����[+"ҭ� (�
��ajf����r��ګ�إ@�ځ��T*������d?r� ��Nt�[U��"����C>C\��L��Y_=�ptQݗ�eЪ�[�
���:��l��[��<I�-4������,�:�;a�W�x���x';2A:d���09�	PT!k����T]��&��$� �?�<:���7�8�ک���6?��2�#���ES�/����5�k#e��];w�� ӑS�h����Wd�����<��u��:�yt+??����j�����t6b�5�� %�$0���x!�a�O"~��k^Q��j�%ٺ1�������)� .��Ǐ���g����:��r�F�s��d ��E&%m<��iql��V���/Rn�ğ)�B��FZ�*�����'y�N�U����Pc'K�spT��.ZƂٷ>=K�K�Ka䡫
=��I����CV~�4�
:��E=꛵C�#�f���'s��Q��P���ty;�%�ԛ�6����� Rlͳ���un���P�یx<~vUO�hZZ}뫓����)�e��8��M7�}�|�E�S[�����	42�� ��򭦄W���6'�RZF��̓)0�9ҡ&gP�6��?;��I�=ʥ@�Ʌ�S������%e7 �1m�c�V2�����G2�� ���̝���2IH
����̈�T$���,|$��G�y��='����C�$�yT-+�8dE�UF�܄Q5A�ֶ��X�Z���	o��wfW���sP��g8n�CI�,�DyV�i;V����k7n��%�H���EB6�Y��̙�kE���������� 1z�/����Xc0�<[̼�����dJ���	���q�^��jb�hJ�[֧21:���ڃ[1��jVonc����M$��A#���$Q���mp����W�n F����n����=`�e7�|g�:ۂ�������y���x��Űz���s� 	5(�d��y.8q� Td�%�8�t���}�T��W��UTT ��eff6�ã��W���HÅ (G{z��� �}�i�L��ɕ+/^�H��v��~���	^�m� �Mo����[�����<��2
�kG�s�G��iy�� #Ҟ\��T|�F�2@���S�13�Z�VZj�l9�����ya��|+��0^�n�I�y_&Y]\\��я1���~=�G�b�(]]^pC�F����l���?�!�4UC$o�xjPZ������N�w��r 	����d�djNN���v� ����:w�X��ٟ����T���G��3�L�{��J�H��uXm��G���V&m�O����B�9zR��,���?�]������(#��]r��n�-�V�}��:�!~���fr:�,���`>��4����8)i2�Bu󘕆�o��Y��Gɻ\9-x;���#Qj�0V���ham{`{Gǝ���)(�OOOZ'D�C~'�]߷�٦Rq��O��e�p��0[Ȥ`T�K\���9�� /�p�j�W))����K8*y�V�(�t��5���5�����/o%����6l�[ ���ȏ�Թ�2H�_w�;�LM�G��.X[�T��0W�j��u�*�h��+�XYQtW��Uj`2����E����@��[�M��j��i����?R=w.�?�x�˩)�f����Ic�k�.��s8*LRy�$�m�ޫ�H�~��8#��߱���ׯ�+�����ǭ�q��5�������,�<�S��5#3�d��̞���!�޹S�N��'~�t3���Y��2�����uq��J�,#�s׶4���]:q�D�ZW�J���toy3Ԝ��ߠ���1�PZ͈EI��0"r��-?���L7�_<�������J��/�vP�d!@�q�D��"D��9���<g�����U��]�1Ӣ�?��5㮍|����zO ��A[��,tW��i~��?
��8F�{�}���ȸdm�t�I���
]2K���g�x���R�S�+[�к�d$���r`�0����{�E1�I{x=��b�E˫�]�.rJ�W��rB�hok{{�d~�d��(
�9:�^*2�<$znv��u�C�szQ���K��	(m��ã�h�� ��.n�S��_�t��khx����u�P��" �ko�B3i�O"�˼٣�2��R�H�Ѵɻ��`��v���|YZ\]*���<�ӷm�[~���0�vf��V�"���֠6��Q~%:�*)q�z� y��]��u��̼L�pe��z�X7'� /��E����#.G絠�P��'D����0I\S �4<?B�J�TRP�K�������F(��5^�tY�����|�m��/�_O�P�TR�0�ͼ/�������cq�HkE�Z���z/���T(�5��'�4�]���޿q���Ƿ0u�!ވu%��V�ʬ����"�D�S���q�K�J��]a���]~8ܼ��(22���w۶n�oj�lR�'����9�=��އ�y|Pt?mN,%A���V3nm6�ҧ���� [���O�Z'�2���j�r2.��lkk�joo�'p�G�E@W�6?"�y��Z�F%~�7 :��!�����ф��I"US�h��0�t�wX��T$It�	��s�Nt�dbb
�ˢ�L珁����8B��@�Ώ��H���EFFƊv,� ���Js�ː/Z5c��Y�
j32���.%*���#���_/E|�"
����*��33�3�nRG�|8N����V��Ĩ(�ߡ�ӛ�u����׊E��w5A���K�VI�{�:�|F��������rH��Y��D�L&$�C�rJ���;��X<^������� �_�5.�z��S<���Uh���y����ge�N_�.�}���d����JC f��8�VV����*�z�E��Z�f��[�?'dG����WRS�dr�?kֳe�H�э�t�B� ��C�E@�Vg
���l��^�"[D��-�#��#�7��
"+YOWIiIA\.��l�6�n^R�G ��"�{���S��Cm��a�ho$����Uc�=��j���d^'o'�'!J������Ĉw܅�r7�9A�D��Ob��7�S��b�r�`�!����߄�����*u�B�-X��<����[3��_�p$A�-���%���T����߿�wm�N4R�P��̽%�T:u�X!�Z(���4�}D|�0�����[��I�3���n���g����؜ȁ<"��&���������v��0�k�{�؛kt+���L�O%�-6 �n��v��MD�$��+�=2��\n�<�XeS(�(Z\\�Gy����)�$pӤڑ���/lI��&tD�"����7����tGv�/��!��-'��?��ӕr�.񗾾~o��0=&c��>ܔ�:l�8�N�8Jb��L��H���;;�3wU�t�p���,��L�q�c2��b�*'3�Tme�?��o�F*�����~b��|t���׬�	]��~����\]�}�zK�W�Nxj�ߣ�O#����e���������t�>�*�:���pi���į�`�j��w+�>�l�y���=_�-s�n	{��N�'���p�������=(�rIA�
��wT�v��K�<ʀu��P�e��ߌ�0�����Ţ���nAgG3+�!�R>���A��g�!J��Dhz|�����S7d�|��,�)+{.���G�*�+���u��9���L�g�X-�"H30�(}at��K|d�����9�M��{˥�:k�/8��2s�T|l�?��V����]��������8+]- P�4��*bӕ�5P���Twz�]S��X����a�s���"��G�����|H�2]�b<j��$sJ�u����
rV������_�
�i��������Gި���׸ty+���7f��C�ִ d�ݩTѽ�#5�S{��o���IX?��ԖJ
5�'L���O#�,�Mܿn�S1i;�ѭ]f�!Wݖ�>����7,�gr/��y���T4{����"��B7����D�rI�#i)V^Ia����Leӽ ��թb�	!|F�1IB>)b#ǚG�6_����g;~�|B��4y7�E�~L6��R�󱉒���Ns��ň
w��c���}��N���8��Na���b����.�_\	R�O�KDߦ��,p��Ɵ�lM@�Ո*0��EDD��H�6��6����8r��zP:""�|am��V�`�׎C�{��8�f��jok�{�����W뎃�{5)���!ؕ��Ʉ��b+r2F:���R�Vzt�ܼh���R�9�{e�dEy�`�ϭ�m���t�Z�����p��a�ӧ(ss�,@l��Lw9%%;}4k�+�9�Wi8� ���XsT5y75o	#�y�Y����}F��r<y�$"�冇�����_�b�M?0����-�k%����6Z�v��c�_&�	%��P�Ge?H�68(��ݱ�9���R�l���ދ%����⛶�M�.����]n�o0d����+���S]S��V�P۰��\�Z��8���vF:0�7Bm�Z�d9�U�VY��c6�\|܇Q�a��T�O����^�L�,��.F��S��z�q
vA�����].�,^iwo�ڥ毎?/�Q$��7�R�G���9��y���P�8�����[1��^I���۸�3��LKRR�w��f��fs���x���5�~��OcgD��3�r����۷�.xe��ҽ����hr���۷�>�����-��d�{��P�ڑi���x�b��9:b�i>׸o�ԕ�/}���h�v�{�e��wiS�Έ�w��e>;s�y }��@V�C�ܮq��M�B$�����9��K㓲�'��Z5mt7�Ȱ�D��p�]�'�{��e�v���A�Сsm�;hf� 5�(X"N��U^ /����C�ꃈ� :o��=rFH��w�5��^챍��$H�$���L��u��������'1� ��A�����
�l�l7�%�~i򓄄���e�e&�����O\��i����pllR���r������亽܈�N���}m��4:z���;vިʋߒ�_etc�#
I��$!Gl6�3/ڇ�M'�|\?z$���h��[�������9R���e5+�k�`i���!���_Z���4��S��8i&�ӟ ($D
�Ç�y�EOE5���ngMh�1�0��*�H�+��40�',A���k��7/K/�CF�իW7QʊH�~�����,��4k}��ݻ�NMCc������e{D��9R� n��c̛�N�#G��]�V��/(,,����s�M,����i�X4�lиGg����B���!UA�5v���Bcjj�:t�/w��y�(�Y_;d)�|c��޽����AHH���yO+�&��ą�KBZ�х�� ����b�Y}Nl#������8A�O��!��v+�V��zU?]���]���q�QQQ�PZ.+�����;�<�}Sa$)-ݶ���- *��+��02giɓzO,�(�<�����c5d�����Tf�SoU�>��^;�JII}��L_ ������kjv��:L�Y���z�{{�SC�=oĈy7Դ(]�4��)�`��ꊐ=�+K�0f�~+�bW�߾HF���GP���5��q`�)ZC�dΝ��ՠ��U�aE����E
D���> �����i~P�a�^9n7E��qT�2F�����%�G�86�V@lKj�A�:���w;V�����Q���j&�NƷf�ut����v� ����Q�ƌ�o}Dqpp��C��MǸ��@�9!#��&@gWWR(�r.>���fkM��b�y� ]"ȿ�P��?��oɉ��n��5���I.Q��y�e���7��
E�8&f~?2n4/�=F�5.,�]�8Ti�4�kj��������H��߻wo
�"��x������������ʪ���b�̢w����qjx���w��.NT�~N���tD��+1�����c���I)*����S��xl|��c�;͠��duy�;��kUP{���i*��-��W��~H &�\��H����'N�Rsqy��� �7��Z����B��4���^�t���F��0�[����ȏ��r��t |�'m������[O�"E���E*����(!-��\�n��+r�Y�!�|�.�SVV������w���m�,j	�g�qp�hA� �*��t����ƫB�`�Ksss� K�.`0������`c�/+ڑ#�V�����)	p�����'�j\d��X�KKϲF�"a|�t���Φ�G<&�
ZJ{z��I�N&�OCC�3�!{�����$��t���\$ާ+(�/��cs����g�!	$a�Q���22n	=�NM�X�g�؋��E`�
��כq��������PkcE!��<����b}t���!,A���k�ܹ3�'����	�S,�����'���<9��b��ǧN�jjj	8����a'�Y���{��in��E] ��-�L��:���#�-��"}��m��OZ}�W��VQjLJ����ϥ;����e�r�Kum�:p]HS�\�VE,���h��(��vgΛ�w t(������k���Y@
����H��!Kx-�:4G{$P+��3�,��ߟ� E�n+�H̯
ڣ�i�0a���DD*�����DB�"��~�����@&j��}���Qd��o޼y2,�Ғ,����/e�ŕJ�};����
�!)����dv4l�Q��>x��_a
����$eV�/��\��b���jԃ�Й��Z��tj�}
|�����zIU�Ȑ�E�?^�J�<8�OFVE��
0��{�וR�������y��%�7��{���e���K��%O�%F(�?9y�ٗ)Co+�WUޕ��&�tkC���/�jb�'. 0��@8A�f9)#���S�S�("0.�k�HKN>���M���n!((�+��߂���횶vF�5�8���Y ��{Q����4w�ǚx^J�]�����?�ܤ���o.�L�����2�`)$ pB����y)i������������N��r4��x5X
Z�٣ȫ(�T)��em..��c��6�>���O;>�u-�SّR��p�o���!ix;����ֶ�~ z�I(I�O,�!>�����WcD�@q���O��"ty�����g�n������U�[�˗�1b��g��Y��Б��Mr�֊{�1/^�O�p!��؊U\_����yd��c�������3�?�"�L)�s�������ove�[˂���g���R��s����GFG�>2G�9y��,��8�u6vv���aV�������fl��o�`	������_D�N������USq��C�bb1#�^����
.�z��`mc��|}-��4
&4>��$���̢Xĝ�<�� ��8�&�}hp�W{����U[;;;��V��B�Z�K����\�.S	m؀�"m���Oq5?�uZ��u��^ּ��4�k�F��*>�VA��GC\rqqዾ�<yO+d�r?�_�JQ��1t(�s\���*�,�W*�gϞ\~�(3��,s{��LW����9I\Lw�7nF�o)�t���_�PL�E�m**ߚ�|!���̋#����3��Yh 3�|�0 Flg�5�7�wre���DZN�f�n�t�B@I�̾�%~���5�;:�~{J�;w�w��λL�;O~,ZM����c�:{h�X��ė��� ���sʆ4��	@�R����8�<	��C�U-,RVF��2��JY�\%�.:;�_��iЭX�qICc_���M=.��g��`=|��CjzzÃ�"ŧ�{Q��}�'}���Z�����������	]ho7����o�m���hvm}m5!g�j��ٸ�z_n�q��/�!L���l�;uq�y����G8�\&�Ŷ���R��U��N�ɜ��x�?u�\9��X�5�n�Ժ�sQ���Z�L���U���ڭ�"��O�KN�,j��9������?��.I�z������6<�����9Y�`R�����O���64I���vmxc^VXX8	zh��L�Wg�H-�j2�-����!5�%���G�0�������d� 4���5�k���5��~o6��퐼�{�\�a�4C���NL�Q�5`cM�gy#>��h%���B�U�a憎�ܥ��;��3u���B�r.,�`��/vNc��*:���[�1����g�e�:�B�-��W#��La�l�փ�е��*e�K��X(�YD1�Y߻x}w��6�'Q4�p c�H��/�w�o��f�?��c��)��W��Xm<ӧx��4��]���mjI�B
���ĴN1���w�@C��4r�znPZZz8��w��ho$�Ы���P�b��C�/W�~+ME����毎����j�\�����t/��Ǚ�N��}e��C�_���LJNV�I��~�,��� �������u;j�<�t|ˡ��8�-��. ����i�_��y�jj>&9ď�2T�!8,|��Dk3r�̋/�vl�N��hD�9��x�ۻ�����OmB��e�r�tu�6�E�u?���xP ���wy$�.׹eWhj���>dNs�;�c����Nq���W�z��� o�>�����]����4X�֣`J��]���T��ϖ�֝����œ����.�_��̀3��u���h^�MJW�9�������_�.�� pw��𓗑w��WI�-746�&y7�O��9�O�C'ΫU��8�����fh|��6C�4�i���8N2�j�K��J����u+�{�߲�H�guh��ДC~�����ŚC.���qMO�
hU�_ޘ�)�]�3^���'��:cù�L ��&�h�c��+ĕ�F�pJ]E\Ԓk��S*RՒ��V^n�,E�4�K�����Y|�	fY�`��+W��o�" 
���JYfa���!���G�(<?��u�~[l�N9ԟ�n�xy����!j��&�"��MO?�]�W1C��[�$���>K�f/�����AJy[hߓ�w4	�!�K�h^Gq�� #��O5�����c	�:�G��s�[����xYzv�'"��7-,���\�`�H{��� t�����e�};m��ݸ��{Q���"���v��w{�RՀ��@��gfBzz�E;�h�*^��7�}e��4��#<^y��4d����V�Ϥ��X.� �������k�3J��Ϥl}nȝ|e�E�Y|nY|�0ڍ���'��{������������N��f�.#Me�@J��-�͑��W�k�r�^ig4�
6�4�U��d�C���F����%�ѓ ����%e�ͧ����Ҝ�E�'�����P!����.A��������`��ꢺ�I� ��"	�����������cp�g�l$��+R]@~Ǩ�4�D�����m�yOd]�����L���E�a��XlJ�<h�=)�m�,��y�y�<R@�0/Y�����G��6�rR��'��>���`�7�K����E��$t�H頍f--ynl-��_�Ԍn�m��|�ʹO(ɛ�@������U���+�G���Z��Q�h��/�s/����]��JJ��~�mcG��y乶}=��?_�S/S>�{#��ٶދ+((��k?�D��q�G���sR-^�BڮX{��Y�Ssaۂ0'�[�F�_�st�};��%�9��"
�j|n�@������iv�-����$5<����x����7{� ��q�F�r�:�=�x�V���j�V��zZ�]��c���]�H��J��"C��щ���8;�1AV�,�.F���7����!4��I�����e�#"�b��sd�
~zz��J�@8������
��&s��O�yN�P��}��ۛ�}������/�N��,�^S�y�r�����}�ۑ����I3�=��e(�P���O�۬�1W�˗�'�"4/8!�~D�/_���Vde�on�zRl
�dI� f�o�v��؉�V=���G29X��ZG ?`�@�k��.�y����l������E�$�:�����e*Ѫ����_��͆o��U���L��=�������� Vz}�N�ɦWf��	N|�h��N����ݓ���6�¡f�5���ڐ�`mD㻻۫��>�#��Mrs�sp�;$���^+o:kh|܏<w���BDH+��ɫ
�2��ow�s��'���222ttu�41$2$���a�1�K�m��\WJu��>y򤐏���sήx,=U�\�S���u�E-��
Y?��`��mpx�}���������r}�D�*�?}�d�9.7Y�^�=��u)��9�����!�D�k~�������5�q���g�5���H��<�P���I硺03�__ ?Nٌ�֫����?��x[:q_l�/�>��Y���n��gF�M###s(-��bO.�dQ���~uq�W��"x]W7h��T�A>��B,{q�ܹ �>9^"�@�C.b�s���h��r����o}�o���u�s4�bS��N�ss{�����-�哴GE$S�)[&
�!�dm>�F�!0�<ҀN�͛�U�`�s�&�bii�"����*L��c\`�x����j����8�����o����"}}}�3���2_�n�S[�93B,�]�ѷ<��2�_�����H����6� ���S�V�i�p?>y�_�T^����U�"���0N�@s$�?��{�0.Tt��y��Ok�z	�4 U�Tʖ�ɴ���S�:urs�����yJzl�k��C!�̾����9�q�2��Kc^g�
��ȋ��7���s�?�C�=VX��(�� ���/{��m��~��d�'��Ĩ�8ᴴ��+Gg�24⾵Ӷ�0O�||�}��-��)]�v������h2�1`�����F���Ah�|�X��}�wڪ��|��x6�>4����H�Ƽ����@��Y��E�cm�`xz2�}m�̹�ź���S�ϳ�/˯���@����a|΄pg����|ۘ7�ɓoJK��i��K�������0����s%����oIB��=<<�@Bu�G	YA�*�,͆��4]_��h��/�_�Ư��J :5?�@& טY�k7'z��
"���-G?'�9����V��l�L�%��\�04�\XV�,0����w�DXC�XI.�
T`C] �t���ڳ;�]�.�=]��Y
e�	ĒL�I�:)��)l��yG-�����q@��]�����pf����	>v������;/iiM��Ŏ,vi 
���-��+���e�b��/��[P���o���x����B�!b�]���0�Z�p��y���WIۃO��:��	h��O���۬o�Q��(Օ�|Y�}8bW������z�8��@��]�bif�'�xL�N���e;y	R�u�8�����.S�+P�$p�
,�]��A�yIC�(r�f}]�h�,���yL��iCV����AC�ӗ���r���;���i��Ou;�z�\�t��5'��dQ�h��鋃���*Ct��`^���Ni�p\߾{��k�0m�B�ޜ�i��E�\��7o~�����X<��\(�8�xQY~�ԏZ�H�t��3�~��!��r�s�~#����?����%���s�"�.]�Lm��Y�׸�w�a%"�v֗-�(�/6Wy� [1{�����Q����FfA�5?γ�}�6�����d
�Ү���/��Ƹ�ñ�U���A|�G���ɜ>5�|*ÉE��CCC̙99�_�=�s���"g��<ʝ�`K�u3o�i��Խ���Hq4�ˊ_��5������-�黺��U�b�!�v��X�,��i��_O�5׮��^��F���^�oyS��NB	�}��1w����Wo>�.U�o�
�8Sѯ`��[��������-DHSӨ6s�B-R�(D����>H�mSƸ1�܄^XqYKK��6�B��8�?RC��][|/�!�c�d��m�2�$��p��Ȁ��װ�7�~\?_pB�X�d��?�RΪ1F��6�(�F�o(���˺Sy^[\];κhebb�2����Ī-��F�/�c\����;P˅DQ>w�ߧY����_��;#�b	�tz��t��S�ۋ]���oɭ�'Rj�V]�+p������~$9���T�����HR,�*�G�3\d�+~}5G��7���vq���P"gHMK��nd�z$iQ\;8���;+���`�˗�q�.�]h��O%ɲh��w��P	G�ܚ��b��2H�H,ʇ�=42��|O��W1������;y	��L7N/��b��Z��~�����VQ	X��<���v�{�5}�. I�L�B�$�L�#*����7�$���8@�c����)�M@:�5�������|����mʝ���������T�b��a�j��J�-)���@��_�F��7�Y&F���v
���t�)��ĸ��r�)���WL-��- ���{�jy�.�ďX@��\�/~�`�R���f�,K |�[�E� ۟�>H�ծ�����m��$�`: ����X�ȒB��|��^�gϞY��0������jJ���\}T�������(������ҍ	�"�-��e��HJ����t�tw�tw�� ����u��z.�>��޿سgF;��:+�Z�y��~p�7�|i.��~�E��ƿ��qٕo��|r��J*nJ��Iq[;"�{��s�<���*��M������(�@H���D�_�\���	�dk�dv�^G�Z�\؋���:ת�j4F��vMۿ�Yt��K$�ŕ��h���6{�Ĵh�o^��4��1����x�y��&����Ծ�M����⼛�<��δ�+��]�*��7�IF�}.s��4�R�{N̛s� ����`w�+���2%*k��^�ay\�L��:`z&&��$k��8�ͱ����-�~�����{���$N�/_V��8$z˵��,� �X��Nutθ���lw�0:O~n�������n1+?�i9�h��Q=V������B�me�BA��bdxx��p�	d�`ߋข��m�J�~��\�w�q��.jJ��� ��ms��������������<�G�;���QU9t��ݢ����Q�{��$��e���n��w�	�E�\�t�&�p�\��D�Մ����l����8R��j��zC2N�Ć;l�������IH
xV��>S�;���X��d`0j��\v���� ʗ��n�O�n7�LAU��x:k�����i��Re�ot�.�L��B��@�:Q��b��q���CKn\�=�Ac�D	+�v9���4��l
x�U�Vט�$a����t���5	
x_���ǉ6�Mf�Ӵ���3������ߺuKp�"R;g��1
;�i�8�Դ�����a:��`�Y��og_����65��eo�y&���BJJ��$�ኇc�jF|k�a�ϐ��8���3��rW;ށ"H�Ծ#�A����u�E�;w�|��3ߧN���o��	�4lڵ\�	�OL<��U�E)I:ن?������,8HKK{[���!GѡX���љ1j�\�����@���m�q�n��л�Y?Ֆ��:��o��)>YPHH���fB�CK�8���Б����ˆ%=��I�^�X�h>�t������m�lm-�7�J���yo���u&�o����M�y�������<���<.p�5�ß̢��Wf�y��`�ǐo�m`9�p.������D�@��-R���ֈ{H\��إ�Lw4�\�-��d�[ԩ���.5��J�aH!�`_�ĩ�|m�S�r�I�,!!!a���j�O�!�7��kZ�Զ���'Vu��f+�c�
��I�� �ށd�U���z���g#��=�!
Yz؜Scgc�7,l��2[�+~j�!�7JP�m�uc@�!p�z�!���\h���%{f�QT��a۠g�efզ�ׯ_z)�{6�x�,0���BB:w�+��G�����o��h�sj%:R=��M:-�VQ���v�T�-�u���t��A�����ϣ�[z�W�^L�;��w; $n�f\RT��#��',��|q*P�`dQ�r�~WTh�:Ȧ� ��`����a����ʘ�����57b�¬Q�R�t"
5��� B�y�۵�* pr�)�AH�r��s�#:�����t�VdED<E����8����u�vC�̍ݽ$і%]��q$frz�C[Ձ8��E8����ѽ��
Ix��:��O�SĽ-�"�:=�@+����>z$K����z�sT�P�=����?����7���)�W���q��l�3����iii�jeG�<yr�c�=�������د��*S�y�?]Ȼ�e�1ӛ+�Un�؍e���~�~��u�>#1 �ʆ�t��i���qٟ��������}ͳ'$$d,�q7��hD�!|9������&�+���E[�v+Mj_!"�G��G�n���p	k�jk[�0[��#_�J/h*�{t�g�6�M^^��b_n�;J�[$��*= �u,�쯞=^�*j�XH��l��{�E��lV��>K��JX�6�Iq��R���{!@j���dh�y�`�yk�l��-��9G'�q�M��J &y��*q����E9�xI]]ݗS�	���i��850���G}�Ap������Y��k�/�WCX|�=�_�}�"
���,�����y�}~]��,53ߩt}{�<3�Y Ƴ��#t��A���,)t���AG]mlX���û0��t݁y�h�^>��Jy빔��`ɯ3���馦�PYIt� J̏?*�N�s˂%�f;��A�k���Quuu�dBCty����'wsU@� 2d�=x��_g����!W
!�����"���E������X������o/RǨ>ܕ����n��AA4篋�E�@H��χ�E�-�^ۯ���m�o��[.�D������b�f}0Ͽy�w����1�	��S�o��λzno�R.@Sz��K'$$|�
��.[<+���i6^�戳�	K��� xI]`-tuE�#/���J�3r���n�X��"��kSr{��I�ݲh���S/A�.�0�8t�Z�h҂�\�ל�@ ���+�;����>�����
�}�Ǐ�+ʋ|�Wj���B'm1��f�Ny��ո�̕YT�k1Ĳ�AZ�Ha�XrN�/�ς���~��_e�Ҁ8���j$58N���53��Nh��S-�󂘴���sA�z<j�/K�¸i ��ꏇ@���D��� �4�i�����1�����

����� b	�7������5TM�.��e_�+әλ���An�577w����=|���OBs�� �Y���\ϐ5�c�&��#.ct�7�����a��=P�g�cw�:Å�������lb�����!RQ�����;��Z�O1f��F@�e���ht��ۣ��;����~�������"�Y�s����Em9A�S1r��j!2%<�H#�&@L�I<<�6����U[���5����s��F��C����;���(��9����c�>ѡ�%@f�;��k0��!!YLe�'ͫ;�ԩ�wsS$:�܏n������m,dgg��*�Hp��(�I�'y�k+�-�u�fO)���\[��w�6x���N)w�=�.1���ʿ�O��>����o',i�[
(�DWo�r���]�hw���������]$"��}���˭���k=j�t'�v߻rE��'�k�Ĝ9gǖ]щn�{Z��{�x��BŴ�M�^{���׃hG�$�_��|���f��>�����ü�h�� ��X ��=��y�����O�8�@�&�bu����с�>S#�����n�S���A,ӫ��h�E�\�&��S �k���-�a�
ہ�{�W���a�|�S�F G!n�t��.?Rt�����|�F���O�hg|��������eof�wJ��s��[�A��6-���R�Ac��T�k�~j�S00H�� ����"�,��{ ��ƅ������ix��? ���3Eװ��.s<�Ob����Ak�j7�Q4q���8]��|��5�r[/� f��P���� �U�V}B� ^�KRV�����Bz�P	�MF�3�����������>i99!mqQQ/��7��r��[���o[�4Q���d`�-�w_Yo���JУ֨	���`��M�<V>�L��
���'��r!�:~�������ԡ��&:�� 5���˪���-��������������L�x�y������pϝ������G�zċ-��w����^]]]���������Τ�����L�����/0��4��E��\�KU�"?��浪0Z�i��p��
)E[S߿�b��L��=F?n��{�G�K��Ʒ�Ӎ�z#�Ή��.�	1��Q��G���?��R7�|)�A&����h@#�9��+��ཛྷ�Lѝ�_b�*Ĩ�&^<�],���\�vG�R��"��9glL��vQ���&?I���$��AL�7���C�+���R΀�����Ni{�B�z��5�.۬���v������#�i80��m�UQt���Ǐ��N��"t���)H���&ZH�%S>�+�G�w��w�T�����\��ߴ+�y<�$D *�s�2l���^9�����"3���>0+�`C"!$��j�����K>t9��s��Bب+S��qH�B�^���c3��ݑ���2S"�#�߳������@�4�c�����?��R��O.�NK�"��jJ�u66���atAAA��*f��� ~c����yÍ�ˇ:U/�?64LQ|�&E`�0:ח�V;�I��deeU�^����)�6��:u�����^�N�PάA�����5��+� 1+]N�f29���ﮃv�����f�E�*R�������uI�@�޳�4��{IЉ��|�)����C�
���6.]��)i#
�K����R\b��J�S#R��O<-H);Kߞ��lqQ�)�4�S6.�etر��"6��_�t^�Y�m��C��ڬ�H ��9�4�R?���
�,�#�?�w�'ɺ��6�oN)���_�>�؁Z���_v�o�Y����c2]Ml�;�G�C-�Σv�m#��gd�W����O�x�����`�7)*7K�x�]|��L�l	�������,�b�LxCP)��>ˑj3����썩���NQ��O����(�S7M��B��;��~W����бj�!�R8ۥY��$�x���N9 G����ɣo���R��,N�5qX�P�����V鵙N>�B����4`˼�O!���SG5�-u�e	�[q��cЯ]���o�y������(�(��}��2������\�rV��jA�������C�����;�;�,Cn����8���ħ7�,��ׯ��?�#ɸ,*])��6M+�=��Wz��:����V2���xgP[Mm(��ε��}�����1,�g7	}!����? C����#��ͱ�$9�����U��C��E��Ԓ�����&����������Ι�����⵻�.��9�0G���&N����[��堗գ����M�������SE]�H�e*k�~ ]qz��r�]�V��gE��NO�����܇---|	))ʨ��63D��{n#$T�866f��u�r�:^���ޣ$����8YV�YVl�|
�,���ۯH$|�:�(�Zw������8<>�Tw��5���C�H��p��q�NGW������h�[�9�^h�ziwޑ/j�r�ұZ��7����=k��j �ޣ��) �kڿ��F�d�~~��J*4�М������*v��=�^|�2ǰ��I��L$p���!�g�О6@֏T�n5�$ǼH٪�ɸ2�(��wdԯ�{����8K,�NuvʎG�;W��'D+�Ͱ��l]�Ұ?�Af#NX8�O��5N�ڕ�l��8�#�������7O�S覀^3��{���O�6m�Y��N-��`F�������G�k�Zr��s`�A��rZ��O�O�tɷ�/F��W.��[[6AlFa�3���q�0|9u+���-Z(����r��6q���Va!��޳�O��m�|a7�4qħ�f����.>�TM�7��mȸW3��(�O���QI.&>^/~5��[��I���!{����I�E����5���QɃ�qog(`��U,	�W��jѻ���+��g�-f�ϓ7�>������n�h'���oO�����䪕��F�xl�*=I����й����0��>�l��6�j7�RAW�"V��
��Bvz��J3jAgBXL7qx��MJɻ%"u8�Ef������b��UI�(�Ɠ/bZ�9@T�.�<�}�����;��q:�,����/�|�!�h�����T��=R���Vٔ��.�m
�������9���O�tA|�����Y��l�2k7����˹�;���j�W��Y���Td�\o�^���t���Sj�[�X����CF��3�Fd�f�/Kș��S��&>g�tw��؝�,4�uꗑ���d:��a�D���| L����;4YE&��l���P������č�����SV�����~]2V�C�r����UaḶ��5ytS�v�3s%L�o.�u�s�HI��}��jЍ_Ihm}nj���Q�X(��Yrن��K }}}���eV��ܯ�u���w�{y�����^�ǻu��������;�m6~ݺ	)�|U�{p۽�Ұ������"�;��^9�}�ȹ�/�E5�(���0�7��M�rN�1<�2��7�t��C��]2\��D�� �4��_�-{w"���ދ�?k�!�����A--��Dk��w��0��9�抇q˩��e7��6��u�n�h�hˁ��0rX&mko[>ߒ0�/iz���/�Pqص��	�n����ffC�f�'' &R,��
����z̴e�q	\;5�F��\���'��;�������R���\���3�Qߔ0f����)�/Gv�5�b�~���1r�+��/�D��X��m�gӨ�!V4.����.�ё���Ϸ��o�t��%N4c�[5�>u鎪��̕�_n�����C3�<k�e[��� '��m���{fJ����r��ŶbjGR�d��۷�ֺ0����9�ž|uqq1�_Ev(k������d���z��gބ��T�����!�����t�|(���;���b�ݣ�����*P+��%#/��Ub�3-z��v
1�Ą��d����8�~�� I��~����fm�������[|ލ= ����w��J����M^���w��Lr_��H�TT�oN��/����5��S��ᆯ��bk����1k�_V�����֨��C����������pǢ���^*Jʕ�����\�TЃ1�5C�ܙF�@��߶m�����54b�[Z�Z�X��_����1,��T�|ߒ�w8�>�����P�5aA��[#�A��OnUV>Aߝ7Қ$��q�L��?
ZfY�S�i���w�1'���N _��<6;� �&��#�Fd J�Wc?����gϚ��K�|�����!@�s�t�v2���.�$�C$�!XJTB�{Q�F�AH\\FW7�@���t��YO��u�9ԑ�g>�bZ�&���H�|Vu{.f��Aw�f!�E�(��L�����{G��e��S^M�W�Z�x�x���6k�7ANDDD9)&��BI�A�m!i��"������YL���ѣ	t�L��7��[׮�4�B[��8?�x�[��c�`����lr�(�����ժ�*�(oR6C5]]��"� ~R!l�4�����2��4��@/��U��M��cp�q��=�K���	{��=�x��А��=3E���m�/�0&Bs��Y-�c���T�z�mv=t�b�\�&��K�d+>w����01V��Fw'#y�DP4��#�������Ы23��L
�q�B�2�F�zNv=���TW��Kȭ�M3p������{�9�/�Ys�'�+*�Eg�����^ZZ"�t)��ڜ0@���o�V��#��n��G��c7�hk��%��N�u���X� �e�>@����0LE��Z����w]ؘ9������|Q�L�18�}U�c�|�ɴ
r�6#lz���LLL�v�zBXƟWكԻm�9bw`_JD�3�I�f��z�-2˴���śuF�,Z���.1�t��7�C�ߔ�y��7"��_t~��֗��wúg�@W�ʤ��R �+�W<6::�>�aT�3�`6Pd��1�:۳����߼��)��>o�ru�O�Ag�&f
"�a��S11�0��8I;�MLL4¿�}s�΢�<Ŕme��,��\c�9��d��Vܼ�E�z�A��iih��Hz0�V�U �ꬁ8�A7+7y0i?d�ܙ���]7kmm��m�����]�Ŷ=�+41�7�ͥ�	*A�)�qv���}ċ�}`��ϟ;s����{d� ;�~�Cv�Q����t�-۰/mi�4�V.+H�U�jȹ������VJN.hƘ}���|���>'�#_{}�o��\�r�EN��^%k�g躼��d��y˙N� e�������x�Be@�Ǐ�H�J�&o����[zO�m"x�le��lD���C|?��>K6�ثvsq!����e�e���f:?�nB�		K��$�`t�kF*4�M��"�h+�#�?��4����F@�0�d|�fuc�G��.�U�(9���t#V��'�>]�ll2 �<�1G�Q�b���_�t�c��1�\v�o/R�����R`*��nT�P��t-'0�kO���� 9��|��ed��o��F�;8VVUјC�(f�����KjT �:����b�	��|cA�EB����vڗ/�YXYu+?\��BS���O�����o�J�Z�l,��L���n�v� �<߿�f�zu����X�&�#$:�0��&�C�y`�Cxh�]{�.�"�썌��Nڌ�Db�k��O�?��!����A�q=��{��3���5��!��q2���4������RQIE=d��uG����1] %M�����qX��=V�������v���5�մ92]����Acv��1Ϡ�n��ppp��*�+�����a�v��,T����Ң`
�=��M&��<~߇�ݙ:ѣ�/!�{�3��$%?��wF ���R��s�+y�L��8�Ç�-&;B=�T���|�>�5�"?�GE;S�ײ�&� �>w�\���Ͼ���ݱ��5c �8{_c�����Wۦ#7-M
m�ە,�be����Ĩ���m���ʇ*��$+:�c��S�j�M�zF�VK��Yn�����pf!Ǯ�	��}�j�l>�Х|�QR�'V�0�������{�2!�}҅������w�8/��$^��	 ��b��3���tz�cJ��������]޽�Y�h�e	�h<}�N����H��3�� ����i98���^�o.�h��Iz._�EC؋S�N(�i�~����w�����J� ��ö�?�������BN�S�)��y�A��{�| Jm�>����B���0�q��c�?F7=h�k���#�T���
V������X��F�ߞlj��;@�r��=������Q_Skk�+����~��emN��|��i�� ��"/�&-mH.�\G<��ȟ?��@[qqq9�"�)��Mg���D�nMRդK�k������H��|��vD{vz�﹖�mY�7�z F�X[��䙚�β��?P/͉��g���!!��=/�R��W%ϕS�g5�����\��W��5=���6.��yz�]�O�����p��33�,
v�t�r2���O7�����)`h��wb�SOOb�|�̳=��~�.�vc������ɛ�,�k��Z�b6>��E�Ƀ�A:��^�b�5�e������w���zv ��7��oM��z#`B�GrP���b����q������.r��Bc��������-8C��B�Py�.?|P޻w�<�Vނ���;,n��4uk�'0	0�7oݪ�n�'!#��b.%���y	w�nA���+�{z2�U�����������_��g]�p!����~��p�4!!�+n�=M�ByԘ���߿��!�S��f�"�6C�.���aQ��?��4�.f���Jy���ge��Y>��z��&�A���8�{��'ǨÛ�K�3�
#�ۇ"�C�V�i�Ȇ3|�����]�~�C��#��Ds���jH�v >�@Ȣ�NbR����ײ����#����y�S;B �o�$i��<|�0�a�K���
#o��f�9�q]�.��֯���r��(���l��y�Z�s9���鎤����nolK8v~ ��u���lq#G<��f�t��=|HJJJ�z�A_MC��� v4��#ᵳ�65]"_b���1羱�a_?Uօ�AjT_��j�Y�'�YS .��Y3���c��%ӫ�]��~h]\CC�����"e}Nl�4<��|���hrz�<i�gV+;�r�0�7�o!b��k���rN�S���˫�:@1J�>��� ��[���Z�����!�9�^ �[uz����ڜ3T�q]+����Jt�e�S,6u/Ş�L�gߔ�����{e�������	�8q��wϱ7B�#�O��J��TTԫ��\9� r���c܂��
�:-S`������:�ۋЊ�>kh�9O���G?�@��y�O���Hv&���E6/�n*O��e���T�����$$	:-qHM�a�KJ��W��&x
�����9a����-&��S����� ��Q ��j������E�����?J�hl�����],�?Ɏu�����`�BS��t!(���4~GW#�kR>��.�.��0@p+>���B��&�$������o/Q�}��\bųdd}�1Ԥ�����2�y2E;�'��u�̫��������ׇ~���߂]n����"nk±��o�����i�~������˫�ys��\�]u�����'�)[[[�a��R�f�^?�]񽲲��?���2� 8�C���_C>q%(L���t�{���{�@rq]�`0�
- j�>�`��;�L�3��G�\�o�#�ᅡr�=�^V�Kѵj��e4�kЕ���Y:��]�;1!A�h�	�4x�6`~��$�t[k��[�n=���a�5����">��@ [lL�e��r�X�-֍��FθFצ{�S!It��3"22�l�
�<���x���������8o����i/@V��5S��6BS���C��8/��������*CT���z�=/��Bۜ��tY�Iכ?��񩈆�N��� ���������ӊ�`��J�(�(�MP���q>|�t]}�ܤXBW7���o?~l��ի)���!/�Ӱ��r2�������Ѓp���v�!�0}�P�En=J��G4�Y���ν���gZ��+(�����Y���B�9�x��H��j�H~No�xI$��}ȓ��	�>��\�����"R22�SI�{>�L���� e��̷�VWW�K=}���-���D$D?�r!�W���Sc��)\R����	����aL^�N�{'�o꽍�v|��T�-&��m�ޑ��!���o-�F�E���0���"��"{[�$4��;��&��j�3����Eb����J+ڗr�@�f�z� ���qT��_�~m����M�_q�Vx�\AFF���E�ǥK��0���������0�2Yk?��q�'h��#=@�Ƥ��6�..�� �����"E�����8&#5r�Q��u`��M����L�q��-�������-S;W��P�l+���f�c�7�����5#�|��q0��@p�{k96���/����@�X/�x��<��1��/_���vA^bտ���#㳿H��=�ʞ*�&椭��+%Ĝ�����k	��/M #�ܞ�|SV^�3000�@}{�3�+�4N����77���}��ԋ�~k�Zգ���˗/3�8������Qw|N?H�����BCA0�9t5zr�ӫ�B��C�M8C��\�v�l���)�G�@����i���j���j~��~���-)��}�vE�[�>��.�Jw~8��i�wH�@o��-����x�Wܰ㔁�!�sș�s�t;�+In3qU,�$�K�8Pl�+ݎ��I�d~+� �g�8�; @�&P��E>� �����X��Zn��3����B�
J���������QQ @�II}��#��{"(�U���R��]�c78.{K>�8.���177wk���認� ����_�%��?l�i��>���\��11?��1�F���"ǵ�-�Y�J-��	�8edA�rJ�NQf?$����7���t9�81=������y�vj�W�<#�ٵ*	10ys��֮�&���;{y��aAhv�潧f�}�h'�\�`.����(�r݌�ׯ��0*�R�>��'�ĵ���n�La���d��Cs��7sB��;��e�ߥ*���y�����U�X�);�~�|���Ғ��Y���c=�:�
��>�[t�qq��`��+z��]tF+?
	g\%�l���{r�=�������u��Ew��}�0w�����]�U�)E�T��6���M�}=Z���#z{C�M�bM�����z#do_�3Z�'��Mƣe���h��]NK**~�d��9��d���Nm|>�O����Z�}�ϋsG*�[$����/�Yf�Tm�!�� $&�6��S9�縿��0�	�+E6���\���4u�,���l-�PN��#����zH ��E^f=�d�MÙ�쪜'�6�:G���ʏV�b��P�g�NA vrȕ"[��������3{���-@��ڄ�_/���Q�n��&>9�,hwq�C�X��G^^&��ꊪ��̌~�\���-F��-�E>*ݓ���ʨ�g�
`cW�?#�zYS���@o�`���{y_���?�(��{�Z[Ay<9����5o؝V��USSSUg5*�c0�k�x`�۾������k�|9v>Þ�n��N��N�ᱼ�<:���+`�� ��p��^��y�N:٬>�+�g��&=�q�~�w�s%$U���\��=F�}���܋��!Ă�V���$�W����8���rj��^��(@����K#���g�\�OmPX�1�\���S�K��F3 �	 ]iJ�
,�ҷǲ���X��a�H�i w�Gj��X��?�q�Nbjjس�ϟ��<�a2��>M��\PP�.�-M] )��x�$�ޯt:� o,?�V������n�^ݓ�1�c֨&<ik�-���6k�->��,:}/��g�br�N��f��SBv��ڭhE�/�R��;��kU�Uu��[9x�<�:�{?��i��t��%��94Ԁ�?��`��WEE�7�w��l�Ll� ���n>�Y�*z]+a��3�ߚ����c!�e��?�7�.Ow�jxP.y_�B�+%�%�ה1Tz��6�g>�o7���%�~ۂ�3������Q{w�|����=��7�6ߣo�XT?��I3�N��_>1h�d��6�~{-N�Je���fՑ��F��gIIkԹ��3���Ï�oMU�2q�E�� A����C�T9��xS�$+�$&&V�vz��%���I����B�ZgT��Xs�	���%�5ҡ:1|�Z�kyd|�M�Z'a|�i�|�d��ǎ�,�����_o���6̲|��d���W�Fo��
'ɤ�������c
&0((AIuM�'�	m�����zteh%!�ya�Pz� �T1�U�P��� 
h6g�p[�0�nפ������ʤ<71I�dw�����3-X��O��.��^�L��*�%O �7��S��Z�TT�8�8]
�&a��d���1l9(��8��c9�@�袓�v�R~��	x=��l�z ��"�c��ɜ���M�k�!W]_�τ��-&��t:a�b����W��l�9� R������i��D�e��.�]ڒ�5���JBLb�W�t8�it�����i/�O�<	O`����SZ�oOS�jɎ�vzõ�.�D1�]���)H�Ʃ�$�W|����@0e�r<6+�?LF��� ��ԝ�t%Ԙl6�c�Gh�akڑOyy��r��~5c�yߕ�OUIE����v�˙W��IC��6M5��j�W���0+<|�f��q�! :̋65�|�9Ş?�S2��C44�1zP*���}�'w�/مl���L4^E�kk_�x�@R�����c_�o4�|�^)�@BZ�
ô����*�ʀ�oIר��N/��+Y1��I���d+�?hq�nFdȚc��X��]_0�zXK*q��&���~���������� 8@`��6���G��1��\JJgw���#��zY�=Й��y�fa��pH��ˮk��~04���qT�t|�!=���>g���`���^֫iiT��u�6�1vu�Q�5����3�F��Q[%R��6~	������/O��] �^��x�+$$��МX�����G�s�"AR`2�O�av�$���]L�/ׅu�(qq\>���W�7�Z��Ł9��>4	ld���#n���ʅ�UUUy;K5`i48�-x�021I=}Z����]Ů�b��䋒��/t�;M^�Qkk�M..������3N�={qө��2J��2��߽��Z�DKv��/rb0�D�TX��/��ho�����]��oI`5������|�3�E��	i�݂��0�r�KKKϟ>�Xn�S	P� yl��Υ���]���:d�9����`�@(C��UZ��c8��u��в��ra��>j�F��U��V?�w���V˅������Қ���޽�]{�ϲ��B�@P�hjv�+`���abZ]/���)��k�Lj�z'!;[����
M6��㨟Z���eO���o0%]�h�a�� ������ˁ��߇Y���&k���01�d��Td���7<�����`jz�sP�u�vm(��|�|�G�M��ƨ9�<ev�I|���ɖ1��3���eee"''�ە.����v�^*)�H�>��y��u���ۊC��y6�{3{8��������æ׿K�z��$&��,ۿc��U߶,��7�@*��{YĄ�F,�bϟ���9��#oa&`H�
��%!��3&��"iL����q�����r-���X�P�B �e(����@�"ۮBW���Ft�m� ;�P����u����
����kq����:��B�:�=#���u9��L9C�%�¸h̽�,]�q�ӧ�n�>��8�Y ���ѯwS-�>�##��n���/��.ށ?�M���t��]@Ω��t��nwƀLF���'Y�C�Fv��c��B�qw5o�^0-x{t/�zo��������]2��0�x(AQg=z���D"'��U�ڈ7o���]�j4P�>���I�3�I��o�
8#Zq���QyO9�]���"ϝ;g���8A���r�N;�A�8l��(6ha����$���L6��(Յ��+��J�߱P`�����zcނ̧��S"�`S�i<�D�?�nF@D��Ny8���nMw�~[����T��:�"P�9:��ϟ���f��GN�݉�復����iK�a@����h(�[=_��  '�`)�32V�w�����)�.n��o��;"�a<���72c"��+���0l�?�M�)C�m�ey��M��W����s��l)R�h���컛?�o¨�r�'��˫L�luU�&�1++���AFL�LO7V���xC8�V a�?YF�h- ���J�x�B�\�jN�^G5�]է�7��1%]������h�ې������D�Ċx�?�}��1.:ҹ��mr���������~xX�Е���D�TeT�洜���se�"�����?��w�N-*RF�6����H�G��T>���0�� J��1�7aJ����j�1@����o��^��+A>
����L2��f]��u��3�"�1T�x@[���F�c�9AdL�5�7��>a���+*~{{
�_WW���f9�����k�lv���,�&J�X�@Z�k]Zq�%w���IT���CK��:# ���IO��U��xbR�����3��˧JpG���[l�8Xc�oG�&9�b��5�1}ή�����>�<�Yz2�I�U��W��'�6t���0���@ ;�2�)7d��m���qbع�Z�nB��j�-�>2����kws	�孪�%����5��������|2'RRR`��vFo�I����zp��o.��~��ll�]�X|ލ{��Qwƛ'��#�)�%@�f�GF��_�4%�%��T	`��k *���k�&��v��?�TAGq?�)\r]�݇�ld�;Ñ�^qT%��\]���r���uoN��� ��{5�����aff�2�	�,��9����=:�c��`F���7�Ο��ucêeQ�BM�se唲���
�5��q1Xz5���eq�(������X�V����;�T6�����[PI)i�ͱ �CS��o���cΐqVzw�~��) �;}��q)V��◢��1���h�X�<AEӡw��Qu\����E�h�S��>�v���{E-*ƨ��L�	�;��N^Ĝ}�`<���>0IУsh-F}�R���ETt���)N��[44�A��[9ur�8'��*	11�TVl`a9�Bњp^�>�:�#����g�0����g0vI���24�g�2D�0ᨵu���y*~�ƥ10~ �a�4��G;��8J\x�O+R�� ��@tc朧�O]��@:ԉ�M�s)Z"c��?�&�! �pqq}c���Z4�abQ5�֭j�'|&SX)�`�1@�>+�ژ�)�=�o������-�������g�+� ����jo+�c���N����$x^ggg`1�k�'j5�)c�[U�ٖ���V� �|}���������|(hT�rŧ���]X0F	o�`"��1ȋ�"S
^^^hi&-WW��X��8��St��8<��NwZ�!B��i���s��(��s[�#����,���򟺖`=�'�3���R>k�s�� .���HFu�56`2�@ZN 0��Ł.���U���L�h�� 1�� 6�����sNE6Q�ϞEA跄��J��{�⅘�#�nH@@p��#_M��i.��2����T62m�p�pG�W,�"��o�k|���!$*������+.���\\t	�κ�~�%	���M<��f26����rˬ/�UKk�$Rp�>�D�k�x
ђ�����ߤF�d8�����p�-������MV�5�bN�-�q�(�yM9������q%����K���-��J�6��*���ƶ������!��$$	nn�Q�t�g��v��l�с�ί����W �ӧO�/J������y�v��lbR�A�4:�K�j�x�A� q�
���^b��;@r��8����!R��0CΓ;N�C������P�����|!�4x������ory��9t6�޽{7��c�������0ڝ���	C�%�����?q�C����m��"�{ ����;
٥�}s-J�F��(AÁ�I[���Z�A)�  2�	{RdLՐq�y�ÕS�On����א��g�^�]��o�?���D�xX��㶂�@�VC���g��-���5t���g�ug�s��tj�|��1�*��)�
t̓�o6'İN ��3֌�r��B���_�0�wqXxKq��ݴ.3��O�]9��|dq����?���w4���Vl��؄̂���^�N��2oֲ�3�R0݅ͮ__��g�.���3Ja))�F������m]�S�q�-�Q?��G���elV&���A����l�:%C��TR� �aԨ&D�n~
Êd@Q���i7^�]�q�K�,��4��˟�� ��w�#;�~����T@>HP&��ER�a�b-*�[JZ����w�cu�顰?]Zro�A+�D#���l�@�V��&�Q�_T5����l�D����?��dE4LZ�~-U
�EL�%u�8ήv����lيs,�^�X��ฝ���1��(ir{j���?]O �o�n��*���`ǀ�p~�E�%xY�:�I������!��WHE�d�H�����+�����Ә0�=����[7�T�N�Κ-j�^M���F��b�z���V��xD��*X� `b3���у�s<������!���0r�&��2��7P^ݜ��ՠ�Ê����R�ʜ�.��N�}�� ��6E���@g�� ��5HK؋��0�X����9�N�Y��RG����i;�z�����X�'	Ө��9����Bt��3� �!!X�6�{4��9�}��t`H���ف�be�U��#oy�:m4<��z4��g��,��į7���vr�/8�`�Ss�מz}:%���B��)Z`��k����ڵGfj�����Eh�����X_�4�A��+�jos|����da>��B�b͸�����4+�Aa��M�nf����jw��kt2<j7��7V�^RC[XXc�gj�®6]�Zf�l���	�f�l�t���ק���K^���C�����՞Z@j���N� �����r���Lj����7�x~��F0�_4����'�Р�<}���G���FI���o�`k}�h[S�c4�(F0�͈��4)@�A�o����Cmq�A�4�S�a��|�.ƶ�v��ƃ�`<�����Rr�����if �[���ؘxЍz3�i���y�I�B��,S�u��wh?��f=�:��*v444�Gm����M���;j��X^M=wvqٺ���ݽy��/��ж�3'2�p }֫����)���1���܀�)���8�~��
����(�>������0�п<���+�Y��M�.T���ؗco!"≚��&��.�-��H�fGߞ��!J�u�i3 ��.�OeUe_c{&��F�wv�)��� �x�ʬ��x�zD��P��_�Iw����`o,��z��uT�E����jPoss3�I�[\3�[׮��c�%/f`kg�!d�[}��5Z���=��
ρZ���ͨ#�5���K��E�?�8�c�U�z)��/��Y�� .��kj�,��tt�U�{0��Ǎ���SiG���R�BN��***� ��w�n,cm���g�1s8m�o=>������dd��hCOp�\�Q|�O���"ݎ����f��Y̕����ޕ�5u-�[��U�Z�,`@AD��,�(hĲ��QE	�@���J�u�TR�%��U��f �[��%�@ț�������{���'ܐ9��9���f�̙�G�j�`���>u���#���˗Q��כt����|
�0B����d��� �{3:z�x����p�`w���B�aFF�m/u��Q�L2�n٩ �ş/T1|��� �!�R?r�05�Bn��F#���0Y�d��g��9��,Y�X���.�T4ڲ��rL۶��eVnIE�������1l�ʓ;}}C����a�v�.hَ�R��p�o��A��;r-�Kzp"^�Ԛ�1��UGk�:��Uj ���U,(��
�P9˩���ASOo
a�/QGk�v����h&���4j���r�.n\=9�ȫ1�u�q�+ 	��D����>0׀.A���W� �Tu?)	e���,/�F��09��
l1��>�����*�m��P��T�EaR��b���'����;����؍�(g.��'ǗO�k��	�5""�.*��	�S2Aɣ�Z � �I�S�Ĭ,ë�7P�.�z�y�X�J�;p�DRǚ�����Tj����%��m���d9�0b`���K������H	�(m{��+���a
"�6�7@�V0p�]w�J:x$�s;�����^;1L��b@���z_0&���=S\�T���`�+��~}i]ޞ`og�����w�yS��?�(��?�������O,��ٓ��\q�ZzNsN$�ơ�n��>��6��lcS@؅�ya��'WU7��;�"��XH��&!!��%h�$(tr!-��ח���b0�R���6��V*h<d�����M���q�el��R8k�����S��ibt,�I����vD[`n˹�7� ��A,�8���x{��`�?��o|d�S,�IիJ��s4i�K�MiPY���u��[���5�̞w������������e=�^A����{���,��\eu�xP�nU\�EFFF8�� �C����i�9�՗_&t�cu�I���B�Oo�XS�_�9��'���!��B��ҭ�we�"Y��U	
<*�R�R����ƺB���OiS))hЩ�F-�}���tk�g�d���~����ǌiow�A"��~LEE�����&��dQϪ��<@8�ɻ{`D����Z�5���Yb.��(�u�nғ	y�P4�Qkk���\Lv^FY�h���g�A��}����n(�i25	�c�Fj ��"�8��"o�@�k�6�ڼ���O��o���N(^��12Ŧ�}1 ��-#k*1
���3�=8Ҟ6�.B1/����L*\��&����?^�R�lHƚ���^G��#%֥�z���>;�V�o�y�ui��$����Q呾2�MA#T�ڧ��Т�k�?���_?~���g�Ș�\�����m�2�;�	��P���K��IjlJ1A�som^�9�5ľ���k����@��Mks�����y Hd�~��4���QzM��K���c�>jn�: 9�<���we%tq����Ͼ��+ 6w�G{x�oJaJU����Nk��D(��Y;��jc���[���I���\jA�X�=j���w�;�|�����t ��;	�4��1�o�U������q)��[\aEY�G7S�-^��<�0l{ɳŅX�V13�C^�<&��w��Uk`�0���~E;�"��F��><�������<~,�s �3Op=����b_V�.5v�f�vRo^[<�itHd�/���*�_�e�h�YE�6Q\�|�^I�R�ֽ��3ؠ�>]�
`.�W}1N�٨��;�4tg�"�1�;�z���e��{����P$V_?GBA;��Դ����=�z��k���*�~�m��e:5�t���O>L��upw*Ʈ�WB�����$4	pm\�լ�^#ŗ��f�)��f���S�(�M.���Ӡ�߉�[Z�r�xG�w���;���3O�i�Y�����K��]��u�w�Y�7�c�#��r�X]v�!����C�w�h� WdS�4���A�-��`T�';:J>�W������m�A%�^|@ި�n�g_����fNY��^�-�xy
ѧ�$��Rmm=�z���� ��Ͻ����T��p�d�&��B�S�W�D�B����0�Ca����0x�SG����О�E[�6P���ѩC������ S�=��`��-X��`_[(���m���
˹\{N�7����4.�[g����/�1D�z��ؙ���9�u,n���m0��������8o ��K:k�7?}�i���2��?Er�V����wT`���B�����62pR�\$;��į�����i4ư��"��A��|��ja3�ܸ�y��,��8�Lv�͍d^��RQ��T&��zL+t�Q5|����o�ս�8!��m���̉���۫������qd3^�=5��;M���o����8�3���ߙ#�x����J�ĩ
��#����]�^򧕵&��n�ΙN�a�z��Y.�rb`آm� aC=>2_�rc�G:��w�"URω��*�I�@J6|@1L��b#��Þ�O��Š��Rf<#���`6��"�ӕԷd�+�$���èQ0V����|ڤB\��V��
f?+p��v����/�8=w�n��"��]��B��!®�d#�`:�+-e��FZ&��`v��6W||����)��@��EVJ5�R����x�ӂ\{Ir�i��ɓ/�G��0�4��7���l���ޗ\���8NNN�n�v��Zo���N|�3g<�N3XWu����γB�cVff�����K�>��ǚ�%����>-�osQN('��	�rB9��PN('��	�rB9�H8X�y�|��6���go�)�����ˣ����w�p�2�љ�����>�7�M���B������?0���C3Ev�u��f���r�@o���A=�$hd���E����������f���]�t�����ak������PK   ���X�j�� 7q /   images/3afa6c98-60d7-4a37-9aec-be07fd386e0e.pngT|	8����R�$tN��J��%������&���-J�"KB�}(�JY��6c�!��G�I��g����*�5��y��~��}?zz[_���&&&6�׍��X?01�9||'�F_|:�����a�t����_�7-���>R��ku41�<�y�������=����%GW����������U&&!&��&���Kָ�ލ�)�N�>,ie�8z�ｰ�Q�>k���]��cr�c���e�kw1Cο�n�r�<��oL���G?[p��?t���7F��J ���}��)�u�������T���%�RtHQI�Ly��G"ovf�}��-��4(pTr�}�һYH�j$�A]�`��eE;�	��݅'�b%�ĦF�lt/�DP�����d�����sՍ�s���-�����/y �ȻX��e�g�П>�J��=H�m,T�k��kT]�t�K�H�`����k��R3�2�Y��O_�{��X��&�T���]U��+�^v�����sq0��96]�D�,潕�d ����6h�8��Z����-1�r���vsѱ��b0彄c�@��)��|�,Q����:��0�����o�t-O?�1�rͮĤ^h����#���M���@�g�p�F�(�J����pd��k=r��{ �zq��-MN[�]E�>Ò��!{��y,��3<��i8^j	G)�P���ʉ!!��[W�JՖ��N�����b���4|���N���.kK��t'w���$-���##��0ֽo��A�k��K�^/�u�w',T��}�E�	�i	��O� {���+m���.�����bmic��w��1��c+ۋay��؜=��H����:�޽[Y�^ȥ ����m�m�%{B��|F��=\��뚞vW[���.��h����?}n���ג+�KE��[l@ af� ��2_���X2�	�n����O�~����Ql���)v'A;1��7�}�Q&��&��#�d�^J�%�wxϩ�"Co���^3��ٮc�$�4b�K���#���e��ʴ�'z����f����7��f.o)��4�;�%]�'H��ĳXRˮ4�������3�q�H"��H�b�þ���BG����;���
��b(�}��De�0$��H��G��j �� ��C�*��X1��D�eE�@���]�,�m��*�$�QB�g�X�g@@���b�q����j�x�˂��ـM��BXep �r�t�ʉI���s�n6H��Xi�"I0��|,#�&��t4�/&wͲ��$�����Ǉ��T�iB�f)s����9�"��'����wB@#1�[�H�=�Ge���y���m��_7�:������ �����A�`a�O�eMS~����&��&^�N쀩ϻ�oʴ�D������$�(�Ѻ�CbC��<�t����G28�H䱹C�xK����� ��	���tw5��D�b<�ˏ����"_a�B� ��B��#�D����ŭ�~�~B�`�@|)�Y��r�L&gIϕw�57	��Z��(F��<W�g?�L���fz���؀g�]P�S��í"Fw�JLF%*R}ߤv�'��L@ri�%|\ǖ�pb�d$�i k�w1�T�Y*�,u*^��v����6C<	b0!ּ�"`K���7��C����Mlh$q��|�@�%6-"�k�OF�&�~�Mԙ]_�0Ҟ�Ԝձ�5���ќ���8vT��d��a%�8�r��3�N�Q\�Z�1:��N�䆸�B*�qx��P����t�@5?��_�0��*9�{R8�q�A����u��E�c�bJ��z�J��D�N�S.t����B�@�/�� �gh�[ [�H�����;R���So''�GqK[���51ӦT�/�����W�*4�k5���_a{H��^�(u��:!
-���Ƴ[
�,��Ä	�~X�aQu�~��p{<��S����*���詎?�A�-}ۯ4}	�S��bJq��pCLJLL�+)財E������[LA��VJ���D�Yb��������ހF{����A{d���������@������_��mQ�C�ԃ2$L��
�FZ��F���~M��q#�ā����׎�7�}�ۨ�ѕ�Q77�����mV�+�ҵqҡ����z��J�Oco�i\�ߐ��{�U�>�l��|��o��!t����������B8v "����>��jF��F]k�\�ʐf�c��1_����ٱ���K��I|���NG��1�JLn��/'�*�ˡ��5�-ڀ0r2={�,��)C����/$��v��^��������ׯ�n��x�����خ���kKۓ�N�Q͙�B��a�˟�CN>�z�Dlh\�C���nJ(Q��������6*:JNV�<g����5�Ԯ�x&�\� J�j�jltۿ��RS[�@"\k���+�Z�]i���GG��i�VG����s�V,a��F%�U˒0Bsl�!���U!;��Ш$����J����e��z�e'$�ܠP�U�Zo��jb��j�|��������9��N<#s������Yt�����B���҃Z�&�!,�(�<uj�c�8���b�ɦ���'���<:::87WXS#�@ԕ���/�?���N�����~jnǽX;f��}���	���Z�*	iދk�}��/w�r�T�����q�q%&JU/�M^��x��u�b\����QфYÄ����n���S鹈Y�Lmm-�P&+mث���x�-h�n/7%�!d(Og�q(v=��E��<AAL�ړ7�L/	v~`rw
~��ؽ
7ӵHaS-z���#�b�C�cw�%
�U�c���!����&�y EnH�GE�=�*�AA�^�sjR ��u\�0p��,E�b�v�-C���������������~�U��B���?ںfDd3��yz�*��k�QY��oPgnk�2o�	�)^k�f���:;�=�����?����	1�����];OI��5x\���������yډ��(�1ٶߔ:����,� �t�Q=|��ufu��a��]�L��/����jj9?~x�%�A��o�q�DL��=��Z�x_W�8'Q�2f	���`I��P����?��8����d#7�A�?nA �x�E���!el�%�4`/�����:�!���uZ���������ٶ�Д������D��z��g�4�l����q�Wf��?��bd�~�?؞�`��!;>В�l�1EX��`㤱��.pr>b�.�3ҵ�w�1���L^�e�h�t/�>����xezi8����KHioo��U�|09̤�T%>p�l�xk��S�#�ѣe�cɴ�6j�5+�����6k1��l!����D[�#+����=��O������C�Ш��}Lk��dMˆ�#�X���q��FN����9�Q��I���k-i�q$���1�s�q��%���2��\�6*�Z��.�%$@=�r޽����x��1_�@#�����..z�P! ��"�q,kD ��
���{��_�q_g�1�����S�@B����ܛ�Ǐ;�ʪ�Wt޸���!
ҧut(��9Kc8e7��3���Z)�f��;v��iK�{�4=�'zY����Kr��6��ntaI��c�y��?��Ib��acK�=z8��x/}^^^K+h��]S/S��7$��iIr�zE��5z����Ծ�h{���ݲZ�gDR��Ӹ1�?U33�3	����J����9���5���[��K$�Or����:�������Ȼ��H�U/�G�h'g�[ ��i�3�!,W�B�ϔ8�"�h4�=�y�c����o�)�F��fb r,��>��F�M�>�V�C�Ղ�"һ��؁��.�����8��9��h�hGק����9ɛ�2␋@�@��|\wղ�9ğH	1��l@e���Je��.~���{��)�2O;��x��n��9uXY����k��ɽ.���#��5�IW�+x!��,IP��߭׬�|�TC��~�-�а=�J/萭��7^�?^VF��F^Ώ�Y@9d@�S80�j[����̇�3H��mi*�Á�氄����/��k�t6�:¦+���k@q3����[R��:�����<=udd@�%I��ef�|DM�ۚ¹�R��TDSSȣ8���'��IR[��E�6�m����0M?����%�^�XX�#Lл<�ƔRP����O;8P��7��������m��t���w�l�^(��X�U�?)V.��@�U�c=ӊޛ��Г�I�e���m���:ꅎ�O����p�ף��*/�mi�tm�w���nsљ��OY�������x����F%��N�tw;� ��B��X8���>��K���j̵��M*Ss����+��%�.B*�3��	NM��E�C������|a������n�����m ߙ
��N���u�X�!ݒE��B���]����cZ1�=.1��jnW$�d�����[Ub��du/��(�"(Ky
�n�d8���ŏ?^���9���R-��fk:�q�Az1`3��6��L�Z��XrLa����r٫W����[� ��D��}}}n��Ds����k����R�4��vn��M>�<@}�6�4�"�~�'�z����/��OK��fwl[;G�X�H �"%5���@��K'q�*�z��K_��"�����3�+����N���*��Ռ�I����m���_��to���e;���M��
ViVV �.!110:��Hd��垆#��GC��X���X���^�/���O`2����Φ����*������D4�=��bDDc�-��ì��m����XjK�]i�}@\��=��O���S*�T-#Qu��(6��K����/ȩ_������Q�xߜ!KLbJ
bw���UW�
�����["��6[���x�!|�0gcs��@�/g���.)}��+^Xp��xbg3�9+�?��b[&&fy�r����9m�{刧�m�X�=���f�N������0����P=qw`�&�7S�GAyoO���9�FءBr#�	ai9*�PYY)86�>Y����N�q�]`���3�g)�c������x�n���R��PD��v��A���܁�>�UI	�� ̀,�Hl-{4|�(�c���lA�b���x�M�k�P������)H,,,�So���9�i�}����ـ
�C�g���a����E����vK�G���Ǿ�@�g�!��HW�R:�x7��� �R��sxb::������k�A�8�Z 
;,�ĂM		���_�/��5���i0�����UF6;�/���qAF����J�`H,TH7\�ۃ��d	�C���sU�T�Wj�R�(5�3d��g`p��c1�?Y�|}���E�@aF*j���NCخa;|r �DR���|.������"7�l]%����V3�l�]�M��\k�9��y�1��#���i)��j�%�\�Ç�pU�P��U0_׫�RW`U���#��{��M�FKWShC��f�H�x�_(Q#u�H�;��_~U�K���\" ���	eZ�\��c���0��ᶺ�3Z�����$:������8	T{�Jo��B��
��^����獋���Rrm�4M4S�h$A����
H�����/O4ѹ.:�����?�2�p��;'	+��@�~zU��5��~�r���#�.b'�A�j�>�>y�-����&^x�S*m�ɫ1�p(ۯ�2�l�3�q�o�Be�y�Q���2��ͩv���rpB�v�Y���[l'P��B�C>�{�St��.�-��!g�c�.	���!����73�OW�UlT���_��ڷ�G�ro���*�t�6V��p㳁�V�����-������_B^�MӬ��#�C#u"B�N-z�!�����w�[�0a�9t�r��l�RD��Pi����?|��g{\��WR$&7לJɣ�ベ~�D���\j��I�Ek�	�����FW����O�*⛮�nHnb��8���^��\J}��A�Cz�=q���	k�6��-x�#k[���MV~�F2��t�p��*>V�Ua4�ܮ���0-0���ߛ���ⳁf��0�p��6�mBl��q75c����M�V�o�X�v��hd@y^�U�;��)ymg��4g"m6��\���q4}u��\�V�Y:���l8q��򄲲rW$;��v1|���O"1���J(f;����ߙ�~6��E���ףX4K"��P���Ļ�d�ݫB��^؏��g�0���4a"1M�`{�`�qD5QO���:/����qqq')b]��u���H͉z�.��]�`o�-���ɲ�$�D��v��0�&O\�<K���FPc�G�C�bQY�e#u��Z�)�xq3�a�nue@<�>q$|�V�����]+-��W��a`���;*� ﶉ=��bY62b���geu���3̣�������+�ŋ�b/9WH��h��_���.�>�i�Z�brk�	{��qs%��3zz�;���˿�8} �d_�M4�����%
G� (���� L-��Ѷo���d��O5��b+�����I��֓�H��Q�B!��]�:1�ߟ����~o$�hs�͟uJ1�Yy&&Wr*Ի��Gr�f��D�Ի�:<����_�s�V��p^'�ב=rm3ǂ�cr	��{5o?�F�p�.r�R�@;YW�s[Wy#�T,}�x`��}*��%r�u����o�BWl}��+���%.y�;�ЫFE�;����N���>`7��z�B���K6���^t���y�Y��,i�s���w�r��A��I29dϖ�2'�50��P���< �$/��9F�xT&&�Y*��f�w(oa�' �oKL4z\���"�Y@C�����kmg��݉��:���bT��y�6X7�k���Vɋ�g�|~N{=�P�}f���Gc%q��@[[�+�C�U�k)�p�� �t���$��{7*1$�Q4��������x���+�|Pz\r�m*�>E>�w��X:�d�7i�3`�%�u�~�!k�^�Y7S7�RVL뒩��%�O~X2S �',Y��j1�*[`%��s�n]E}��5�pJ5��)��J��UBg�D�}q�gOA9��jp/���ID�r^<���F�H��l��'�r��+�&�RĿ�'dU�6&'��Y�\L>���NN��k�5�|�C#|��:�d�dP$1��L`~��<�Y��Q�e�NJ::�?y�U�ci>�<�N�u�tQ]c�l��§�3S��"����{��m�c>��ⓔwḑ��|��G�E�+Ĝ�l���(W��$�O��k��?�9:2��Ë�n��Q���!I���}~>'H:���URG[�\~�_�k�������!�	9.��XY= M	�!1y��x!T�L$7�����؛�>�%�k'&uc�����[%�K�~��ȑP�oT�H����1y����z�����'��eJ�4����Ѣ9��`w���7(�,��
��Y�)����k�Z����̍�-9�U����Hd���+�0 �#���`�0x�?k�4��.��I��u��e;}�d$=��u(��YZ@�_�{��kj�Y_9�� �?��o�D^�<J�V�s,v�l����I����Y�"p���u�G���_g�}��FA)�"p�Bi"�W��aX0P_>�����N}W0��kXrwT�)U��D �Ĵ�Ĥ��Gv����О�
��B:<<���kIz,��r����c錪��+��͆ʞ~��o�i4`S��~c�S�.�fj��^:�P<���<��pn[_k��|�U�K��:�(tؤ���b��	���D��p���{Z�p_��+��Q���Q���u�M�D�#��PW �Ĩ�w \V�D���� �c~\B�RA�R�J�YA
��E
�i�^y?d�⶯���A�oҏ�/�C ��.4c��JM�J_��-2�5&�S��T���퇿�ª84�=D_��ec+!�P#���;Os畁FMP�{�ʼ���hVE&���������+���FF��+�M�[�9��`�k6���cY���[�	�>n�c��G��}�ޘ�H![kW0���Oց/rNV�� )�����̐�֠}�*L_���?-���E�~������y�u5�Ǣ��$N��T���m©I�{K[�B��-0���/���{6����@��%�c�6bB�c���Q_�Y�{,���$��+u�gu<@�gǑ�Y�����c �V\c.��Z�7n���}G[�D�}Y	[�������|5�����Z[Ƌ�\E@}�IY�?@�}s��&F�#�r2�H�U��=!����z��򍓗<Eô�N�\�����.��"���Ȕ{�s��L(7�S���ؠ��?�Ϊ70=�u��#T��ЄWTp^���;��b����c�Y��-��	��̠���h�١-{$��KtS�Te���1��$
��:�"�%==l � �F)����J
}�b��_�]��z$�޷LG[��)�� ���{�Ѿ �����o�=N�b�. uۃ��O�k�Cpp'DiQV}���,����Μ	���PH^�G�e5���4N%&N�eY`�M�� ���8*�� ��'{�c�"��7p��$|ڸ&��2�C�C�l�G%��x\~'a& �ݓ c��ߛ�w�B>���x���bv�9��u�����;�^c$x�om�ɍ(?�5�5�@sUUUy�M��gD
���VZB�)���B4 .}���5�4g<�np@���α�@�7^�m������}��κʘD��2���+�u%�E2���A��bA�M���x&��2m�����A16�[P�����+;�]�Hu��u�}BK�t�9Zm5�$���<Q����@W ��_H�)N`���R�Q���	���A�!��f�/<�Ϥ��GEEɪ\�}�z���d�r�W��x]�ɬP^^8%��@��� ��_�| |�t��)�x�z,�^����,���~=�o8��H$Y�ښ�!H��ޕ���,3�~�(��#.>�r}���O�^�5ꗉ���Rfy����.V���p��k.@����γz�֝>Q��ת��jq�F�C�]1�IɅ�.�#�O��+��C�)ej��gR9���ҒS�/-u�;i>-W��[���~��m��
[��BR�ɨ)]�c���j?��N��/���<��Cl��L �����$~W�t�hеV0yc���,�`��i�� �y\4(����q^A<���᮪[WܰߞI�m��Mx�����S�z�Ma���n����<�h>Ax�٩m]�^΅�x!}��)������tB�>[��o���w�)�o+�l8�@^b����Y#��p8�8tŗ;J=S��C����e����Y9�R�>\���י^$'�S�n뀹Sz�nq%s���XW�S��x���(��|?Sc�V�i
����'�'��4����$|����giNO�-�e����f?b����� �=�q�V�����K�q �D�����!�§/��������g���:;|�^�r�p���d�#�2)|\ܪ?�k�p�0}�x�]���i+Pպa;�j�/�n��ST�q�u�iC����ދW��m<�S�8 ��b��ղ����=�I3���u��kYx'zk�#3.�u�E/S����Ew��xxy1�?�w��y9i��d���[e9�lV4����ւ�SMC���U�,�c	�`,!t�d�ᮧػa	�7�r�zU�vv��פ�������t�@��d	�Q��ge
37�d.&��:��GP�����_���������Y���E
���m�k�;�x�r'MS�kn�Qu��A��^�Ҡ��������_�׎��C�[�z43t׺�BeC�9�����yTܗf�ʱD���iy�qBxo-��{��M����+���(�W�M���FkW����Me�>��e.��1C� 3�#Z-�G�Xt2i�F�%C(!W�EX��#j������OK�ǒ?0�7t������H�Chm9bO7�^��
l���9��n&~�����Ŷ�_w=[T9_Rt��D��	�R^^�rQ2�X��c�E"S�d��_����w�r��r��9B�A��D����6�Ča@���"KE�=���F��0]F�,p�y��f���Eݛ����_1��c֏�" -�)ht���9���\X��e��w���Ӝ>������B�*S9p���
��.GL�<�@��=�ֱ�/ҏ2�DbB��n���V�Fd�������?��F�D-|�`q��x��c
���[ȃ2f�i��]ڗ6JNK�]�[|��viuB9pj��)88�21L|L���<U!C}U��Ω���~DI�
9�JZ敻�nk"?i�u�.�k��z�����^ʞ��l*�`�qm/��LK �����7�߄�?{�������������O;��b<����.?@ �^��P' k�ڹ�zF�4j��A4oЏ�t��RZW���!Сx���I�XЬ��,������K����ʆ�7zՋ�V;`{�A� �ݜl?R���H�_f����ـ�2�X�зH֓[��n��6��ϸn ��u��S0�c�WU0��)�n�'E,��]��]W�h��6�;�zh��dT�������,�C��e���lޑS7TBˈ�O�H�g(��j�r�d�?>����r���'���>&�Xi���ݱ@1���o��,*3�ѕl*���G��������p�{�Bd����5��9$	�|!s�u�VU�03�n��|�}�D�ggI�6�_��e���A=>	2���ze�g����ۤ͝����/rS�M��$���V]Y��;ԡviu�:M{^�k�Lc��a��d���1�ßΜ�A'���ڢ�{����$�hB�:�/u���@���� ��O�"}���ݤޒ��|�X��I�ORA敘k�t�^���V�Jo�t�$��Ҭl�L�bA�Jd?���5E�QH���:�����:�Ҝx ��s��øW��ᣔy!���{�U�h��\Z
�O�����OR�����h�,(p���v>S�O�����8z�pU�����hW����B��C9�"�I�w��3\W3��v[�Q���NM��yv���#:LC}�w��v�m��o8�bMB|��+\�e�̲�IS�?
�mZ�� vOf�&��Hj��-=G]���RQݣD�*v�]m�h;�]�IT�;�9�Jt}Lo~����Ӷ|n�z�Hjn��'�<���?�Z���*�wֱ�`����������s��i{�o���Q���9��>�Y$fe�v��������7�_��� *]kL���I_�mh~��k$nk�o��-���@r���o����z�����nb F*�l�S�̘�z����""��	5��5Y��㣣�A������b�]{��9Z|5��=-}&����a������@]����=��M�lt�����{o"������	�+�X�#1Wj�^��KH�P��}���>?!�7�	���f�Ny%Q>F��\@P5{�0?�����ڥ�@�4�d��Y���52�����Zn�;t�7��q�ӯt����x�+��x��kBR�bO�r��p�m��&�j���V���&6��3�,�~��p�OE���@'6�d������˶����έ3zz0�yi99��j�a�\���V�r'2@BR�\&��s?SSS'W׾�9����1����a��
h���)t҅��x{��i�P�؀faW>�^E���[��3��0���;�)�8�o�~7�O��о �|
�����x�l���,g�����P�|�i� �i�u�wR�X�A���!�D������Uν!�G[94_np�@ y�|���0�\5�����Xh���D�܃�uW
]U�߾e�͑�Fp��N���k>O(�y�~-(��ƹ��q���c��i:��#����&�sE~�Ĉz"oP�S��q�Z`m�ͱ�����������"� X.,��Դ`.����j8��Z%.���^�����m�,��\R��X�؝�B������NV���͝O�$U޳�����4��W�83��_ۊ܎�<����ӽ1�#'ǑJ2>Z��<�-����|j��<jG��ER1~C���ڔ�m�Z��>ɂ�[�pQv�1�e�D���Y'W�N��&�_�rq��]Q��u���O?�?�a��/�rlt��
�0��k��z�+Es��
���!JI�A�	���c��qrjj3���n<�@/�==8H_)��&�p�&�V�&��r�������F�
��k�v
�pB��T� �� ӊ��VYxdhp0Yr#������4�����]a�����
LqIIߋ���ѯ��uzKAΜV�j��
�I�����w��9M�
S�$S�,��_1�t.S'������T�֐�^�z������	����������+�[ih��Պ0��j6��2����D��!PM�����g��YS���EXZ�������'�5����gh�,�{�|Ҁ�xW�^��4孤����D_٬�Ԣ{�n
��^zNkZ�ƫf�/RBqY��/�/c�h��z��v�tW�������Q���WRZZ��V�0�ox�����E�֪�a��^�����\Ta�V�G>��Ê��YDݶ�7�U�f����..�箮
���7��j�s��k�z����, w5KNV��4a�l���蓶�'4�1oŻ>T����� ����Q_..Z��?R��{�SsϋSs����TيV�����'�@`��rd��D�\�����S�V�+���2s9U��x��(�����F鹽n/�A��!:FfZ6��s��q�g/*�a��������;(������H�ڔ��F*)5�х&�E{���ZYZ�#�g�_e}���Њ��R�����&{��\F%��z��J9��ck\||}:^@D%F��p��[Ѐ���Hs�����Q��n�ȣ��ô�5���q>���[)�R�#u+/e�q��Dt�>v�Xz���F�}	n���hɴi#,��Ʋy9��C���?�ySW�7�57���1����3�� �<	Xk6���hA0ƇE��DZ��3�0#O� ~Q�8=�_�bt�>�v�ADMM��+Ǟ�[K?�۵���UD� ��9H�k�W}����(���Y�ؠ�����	Y��~z�Y��\�*��"���jԡL#@�;��G�'uΣ�3�S���U������L,,^���a�J��� �����<~|��TS���VF�ݘo�G�ƚ�z���jߣ�	��M`��Z���DJ;��S���+(�U���ߚ9��My#u 1�G���))��UTT���t�X���}��_E��x> �<f�͇of��[���ײ�Fge[| vD$F�'������R��hv�De �u�x�j���j�j�:�boP�.ij��ϴv�B�E�)S�����{L��b?��x�GM+Ԃн�V"�੹{+A�����"�9�Xi�W~�������Z���9e��2@"@�9=��B��$2�}�qYÔǣ�.���yV:�ޟx(�d�.
�nM���(ef�Bh����.,�|�g�ں&��#cK���bqu�V�N��\��gqql 2�@'��[J�u�HN..��<<�I�}��Y���U\�F{�K��[��w�T�܃�s��l]I2O�W$D ������τ�Xmd���ˏX�v�M6t)%WD��]�:���� �ޗ��D�J�5�#w��ź�{�j�S���.�ړ���*�&�u,,F����"y��M|�N�`P���8�a��jPq����-(r�Z���Ļ��TaC##��{�]X�|}�0��;ø��� �<���[*�����<�0%��P���:�S��^�;_��������ȲT�Do����V�ogUz�A[RRn��!�hx4�Q�N�β�Zh]��| �X8��C�moz�{���h����k����������#�éiy'33󟫤�H�4U0��޶���P�|�}Krs�,�M��-��T|�b�U�	��B��.֞��Q�!�l���1���T���eJ�v�>��KL��W?�KH8:9�k��dikk@E��%`<�^�-o��@7T���m����έ~N�C�zQ�X��}�N�Z^����8&&�`��u���p%u��ř�}Ch��2[����o�JJ�'�^���7�#����>y�(��U]���X����1���j+xOD�+@��G!C:�����񹦔���"�NN>�W&$q�W�W'�:;���"��9;��Ղ�=��گ8<�Ijp����N��qJ���H��&$o*4�0Etq1���&A��W�ׂ�N���2�N��漇��_W��U�9Sz�ӧ�~.���ލAl_NE��s!3��R�>��|LaQ!g���HХ}�P7�A���`���1KP�\ �����,�j|־�m_�";����C&�0�����}����T´,"������^7.xF#A@m�@����G2%��
��˯�٨�h���=+�W��x �����%���(y�`UxI�E�[�����h�k�R5XYYY\P̮W��������� l��,�~5�{�_��Ƞ��_�ȠJW����x���]��ߙ�lӥ�k5�,!��Ԥw�j��1-fqU-{;����7�o��,R��ŋ��mT�,�f�Wh�M'V5S������\���MRG��95MGP��*�J�-\��ÁޖII��3�{w�Q�oջ�B)��"-99�6��%PC�b�r�2I�@
��|�@s&�G�/���1O�}!uT��(;��jPD`~��[M��g8�u)��?E�X���yg����y�Pٽ�v����A�T�:b}&���A{mmm�Y�i:�����pXk[G����H���`��� g.���[7�yy������gZ///�e=1�T����|���=�K:���mР�Q0����{�5��.+M��-&�@Rw�݉�)�ʄ���w3�d�DvRO5p���th���Uh�d��xys4��M��\>�f��?<\�]��Y�k�P���i��!�����|�}H��S�x�%��_�~y�M0���Ϯx�zp�8�M�7o�� ��L@?�x`�ϠEx N4�I`|��bȫ :%*E�M=�a��Ӷ
'-�dz����@�H?�����Ĭ�]4@�����V�A{��b|Б�jAw���;io0��x��ҷʩ}��ā��I���=-������;+ |ՙp,B����'Yގ� ���hwu�Q+´P�=�����{rRc�C�j�j+M�X�����T�k]`}>DJ�r
Qo�� 4�?O�'�խ9㶴����n�o@��^s�j{�rek�3�*���eJL�@�=ff153K�f�__��d[��1g���ރ��hW<�,��e��0(��^��_�RR��2��bb���������i��^l�XR�0�ｮv�rY�W
���	����xjb�E�����DJs���vM��S�KG`��h�/�5\Qv�j��UQ�s�W/�&s����$��׵h��ۖ1��j-#ݮ�Cn;n���xA�,?>|�I�~Q��q�$B.Rq�|��~���k({�^i|���)dė����h� ��C}�u�dŚ1��fbfZ�=3��~EC`�����P�3��D{H7Qǲ��u�Г�.��Bh��zj��h�o02�4O�3��pGgg��Ӑ�.Ӡ>�sc
`�.����h��ϾރBͯ<�)���A�*��9�'k�<�rm�:�DҀ�q�ݑ�t�pv(+-��r�$m˝<��m�=�{cN�(�f�/��@��wH`�W)�KI���+p}E�Q���r�j�R=�ԤfL]fpF��ݏ��0�_���ms �4���������1V�z��k~�qm��`�Y[g��R���r�t�E5`���K�9,D��*���n5֌ޤ�`ٝ�u�Α Y�=85�3]\]�%�e�����V谬�tE_�kKkk=�\UF��%@b�44hQ�["��Q�����ktx�#]��D��J%������ft���)'u5��+�|�WRRb��w��k���`W���I�fcph~-�����������MM���"�����&���
9���Pq�E-� vܻ@�}�zj������l�+� 3͝+��;)ꚺ���U ��*��C�
�|�d����B����~CqH�mi0�U^__:S?�+P�c#����s@� X(F��>�_O���$�}T������}/������@ې���lK+��#�5�e���)���^`	+�P��>�ޛ��
�S��\̲��Lo���T��iq��)�� ����X��6���"7�a��,��b�R��?�Z�:|ʹ�e��;)Ė;�ַ͑bc#h�|&�|}}��|��¯�b�\b�/Ў9��EL��צl(�ͣꗁҚ�a��B�7�aU���@ �$�/t�4��K:��m�pv�1���0f.5+�]����w��?�{�PTLl�qD��d��� ~.��:��,m��&?]�P�+t*���ҫ���-qҥ������r(�fߪ�x���_�~��9�Ƒ�h��>>���0>�����i���]Ɯ��ۡ{�������LR
����t��JGlV��#v��*������X@;(c�;вK�2��MǬ�5�Tr�07d����.zP����"eTY	���r$��(ϥ���={�U���>0
��C�/6�QaO?8�[�#�I7j��{U,-ο�V�_{.�lLfu�L�q��ʺ�]D�a�[q]������z�t�������au���e�t��+��jVaTM�"�N;��* �5�@���m���� ����I�WB1Z����|cj�)f�i7DN^�\f������+������冄\5�n�n=���I� ܞ���CQ��R��|�	�$G�s��0q�4��L#��qqq�++�^����ј�*���VS���F������gttל��D`�۽H\����N���H�==�C�%$$�Ӳ�l���N�.E"��|�{���.Ćª�o�;Xc���7&�6li���Ӕz@髀#�vpo(r�>�174�p�2��)j83�tt�4�T&<bH�\UY��`�x��@s�_�ퟙ����q�l� *��ފ�����MQa��Q���8�q5K �P�,��\�s�1����;>�q�/��m\��4�W ihh�'W��w���Ѷdic���������]���oK}��˺
�p�%���H�����+ `�ެr����**� ��/�QӃ��*#�1��5+ P��^c��Xh�Z��V(��߾� 겖^�g�_GT,���|}z�fhS��"�ଘƱGޛ�����t�ɋ�PYi��i]墼��|�b�x�2�<=+Km�4r��D$S��8űwZ]��-�����(�!^C��Յ��r�c�[x�j�C17�]�1䴗��m�/ի� b*���O�u�lG�5v'�9�y�����d�rs�?��t�>�Ӳ��oSX5?b���4���Ǐ�6�~���tn/�5k�;1RNkc"v��fKϝ��ȶ٪7K�,=}d�����W��`����^tIq�m[��>>^���b�X7��m5�R�!�yx�������f!;Z;��SWA*���w��/���ŃSX���͎�>~77��70	��x����B�\��7Z�&B����=��J��aT� TTwU�"��D:�T�U�"�UJ@QpE�ҥ)R#-HJ�H�  RB� B������=�9����3�<ϧ�̝��9���V����i
z� rO�X�~f~���p����w�;���acN�I�������l���ٻ��<��H��cd�����o�ÌM}�����]M��h�۷����X,/\�|c�������>�uwF�7nN/-���I��>@K�ֺ�G��`^�20X�? ���<q����o��"��{/��P֍�:�D�,>����j[X�>}�I0	{`e��|����ۡ�*$IX�ms����ݾ�h�����(erwsb��q���%�m���ħ[�:���6��Hľ�H�������$ܗ���&�]QV��ؑ��V�P*p��w��k�r0�ި�?�w��Ӹ7ο��k�-��4�R�5��:��؃��	Q�����V�N�T��U{ͬ��/���#0^c^f�O��~Ak��uy���a����7e�ȯ����XH7a.J�pG�#g\ϐ��(�����6�����O9:;�J�Wp�5iNO�(ݛ,P"�<Q�����[�%<:.��Y~~����m111	��b^~���y�zx���t�&������X��<Y�7��mT]z�a.*Woz�!����:��`�G)��2O����w9�o��t�J9[�]$v������T�ؕ
����(���`T�|��� ��,z�dR��Vu[\�����n�~���Bi�Ww۴��cR�����DcӀ d��%�O-T"���iP#=h��X�G(Ƚ�p*�4ePZDMi
�ˌi�a$��|���9������X"�%�H��I}3��(�]4>nc�u�gfF�>}  (��O�@)�W���OTA[�eWKJ���
�l��1H��_�!lRâfm�ߤ�پPߑ�6WW�Qw=ټ{~^_]C�� [3�y��֖d��o�"��ȧ��	9<|(E5#��Ln،c�$ew�K�:�,{&t�"��Ǜ6S%��4Zk�fY&�W��x�ӡR��!s��Z��hm$5�$n��A�l]���r��3)p
��|���c��7��u��G,�P5�y�8�Y.�����
�<�b��
@{��| ���+G��}���h� E�
W!k1;`�|�w ;���b���O����_�Ii�Fӗf ����h�������Z��%���[�.��嵬����gT���q^cMː��.$��.�k�v�NN�˂��y��<�j!���y�SJ﫨�
Wr�HL���/�n��M���C�E-yy��Z�4��9�/��'!I�J���r7���\!��V��ޮڊ�YX`K;��@��AN�S�r_/����?�1i�!�9ﷷ/�~T�C??U�F�W}T��VE��Ң�`��Hr���JuH^�{�7�[ec4=K%ư!y���!8{{{��R�;��O�[�c��@.)Oe���{^��fL�I�a��U�&#Eރv3@�h�!0��ɹ��|j���gf"m~[�(�u��S	�9'�h��\d�7T��-�}MH�P]٥�� HBS��d���߂��Fv��?:
�.��rf�K}_.����ގ��xy{;�;Rf�q]�,.�/LT�v@���&�2oqѩ_�{�DE�-|�4楮�jR��h���P�{[w�����I#���Q�*��J��ȍo�7�DiS|���EA�~ve565U�!�1�]V��f����~��2{�Fä,��{<����>B�g��W���v� ��mַE�- ���E�JYȺ �e7����T�.�Tٿ�76.n��#и�mN�!�W럤l��g�y�\Kk��H��|K��wS��2��<�>%.��U����t��p~���J ��յ����70Kg.��ދ4��"0"4��T*�[ӂ��5���0�P��+�R0~s�g˪���8�8��fU�V�p@�.|jM=Y��)N#E*kb"6S�C(ܳ2;w����s��@Y�Cc{����0���HaLt�k�����ꩧ�,HaA� X��_ė���\�IX#��"31��_J��Y�5L.xK�,n7�(��a�\ʮ����0K�������"Wr�Z�����{fU��l��w����D �r��Sp9�����m��V��!^��9�l����OI���4�5��˦���P�����&���d�����_�Z����<G7/TyR����Y�U�ۜ���We��4��(�a������Ll���"�fUQ�E����Ռ#�f�c���w� 1jd��~?(��I�HR��݈��Z��]|P;�kə�.@�I�:��WĀ8ڻ�/��37�N�2#�ڿ����b��$�nD.w,��6�J��;���#s������gf^����{a�
��G]�>�F��X��������}-G2�ʓ叛
~e�� ��#������e!ڴ��I�IL�QBOV뙘�|e/���	�/�jjX�;�qyV���ׯ��)���׼�~���wrh����B3��I�^BCG���19���LP�7'Bڎ��Z0T7W����>C�Z�쵢�N�L�7YG��:��\*9�^ZT�Owe_�4�3`�u������J�d2�Ex�J�T;dw��i.|`�@�����޿ln���d�.uW���t�?R�,,6Nݖ�!�$0��	��d��4f�
���{��-t�*P3V��>��/T��ۛ8�\�pe-��w�F]]�K��K�.9>|hz��u %#�U*���цz�K�
�z��c�ӄ������u,�N1�2����>H3�oG��8��e
MM0h�]�2��������(>�� CL���Ư9n�ŢS�UO��N^ɪ����^����s@��}H�ԗ��KE��{�B�Z詳bs�2���%ҋ�b��3�����\���}��B<��_׍��Ō�g~j��@���&w�hС���(�8�w��w��5L����6ȳtIj�� >>>�����P���paaa^z�v�'�� �)G[?��u"�<��T�H�e`��8�Pݮ?�H��6g��NǢ4c�����2�*Ȟ�۫o���"R�.J�~�%xwh�hHp=H�4N���ʳ����+��W�0v����{��*pL��ϗC�U�2=m�7�嬾��!�K<D�2�韮�
�{�x�H"P�ԥx����(����5�ӡ�ɀ(�@��XX���b��?#6/EC�'����L�&���E02m�����QZ��A&�s��Z�72Ҷ��2%�Kv�tt���SL{=�d%�o��Y��1�{�Ҕ�r�1W�b�k`Z��j� @%-}�H|�ߥx|�u ����������]����������L�A��W��RY�������/�G����,,�.�4�l�6��:��;�7�2���^�]
Hg�?`��m��I��z���bm!n[Ǉ6�"1v��_���#o_�Jn���/��I���՘)�BⰞ+ҩ�>y]���[�
��7>ߘ�n�e7�;b �ꔟ���a��h��I�I���F0ɳI�3�Tt��퟽ v�ֱ@�s����%�����>��v�j��N\�A�$�� G��](?e}��wg�%jcw�3�	'u{���N���@���+��6Y��^��X��ep/��X�Ԫ�E�x�O��V�M��SP14�50ԩ�<">����<{���dE]���}9����-�����`�8ϦDP�I7'���g�0��t#7~́�r��_���P�M	�V 	�ChRQ�7����?�*�I��S�d��쒰
o�U�oF� ջ<Q����uK��(�'�	��4��2Z�ڗV�)�v�Qԅ�������iC���[�f����e`e�-�c���;m�{�[���*	���������)U8DZʰ*�sH�D_9�g�跽~�k~�/�o{���4�/����y��-AYB;qnſ:!њ��q�&�]�c.�h�$�̼�rX�&#mCp�=x��?V5Gmz{/��}~~�Q��������8��X�� 5hc5�������
>7K"&y�6�����n�U��n����Rxe�1�����Ǒc��"���������|�q�x������b��(+ ͫ�a��566u�8���w%Y���7W���q��3�$��>��X{	pߕ����or���,��éd�.�����=0y���&���76�f��-&W'__#]ݨ���R=5TR��d�l���I�����jX1r~�(3%���b��9�,� ���"��Y����n�Z�_�}�N��f��tH��MOgꪶLʮ���*g�a�e�=���}�$P��B@	w�����#�� 	M���<+��/b��CջE�$%F@����CV|{p���ԭ?W� �kt��Z!�`��;x/˿&�R�x�k9������7<g~6:S�O�5h>�vFD�������y/cY�N��0γw[D���_q�:�kCZ���TwS�*�R�d��o[�ޱ(c�j=
��j�2�^<*�hJ�u����1��mm��5�p��H@��6�4[�����a����5���"��G!�Ɲ���6��2�*�
��?��*������o}���iM��%?�x��6�^�V����)�H+�{q�.�v�:�C�����~	�����^���x�UV5+���}:\�:T�9IF�����l�d��|~D��:4�r�ad;�腽`�q��~�(����P])��Ex�=�V��(v�5�~��	�,��f�*_�l�u�L�P�O��@O�� �D�E�t��	�$h?��x�Ω쾤QE�	�������R a\'S&)!g���R.ƒ��ln� b[��i��'��C.���i1�������&��k�W7NPF�
���z�
�TV�Ju9e�w�T��L�#g���ي� �Og��ȭ+�`�'ɏ̀����1�<S�|(~}C�d�~�~bN(��oM_?|�]h���dޱ����tV��x��(�=�_��0(���Ac�j�dJ�7d��]hi�!D��Oٝ'��u~����/g��ů0:�v�*�����"��
E6��;B���v���?*��QwX��)���b+^k����5�w�>�&ppk��_�J�d�*9W�%kP�w�9�?)�A�����b4r&�`�r�����h�!�t.�~[ZUQ
z�N9nv�g�����Y�$"��w�,S����s�$���@��w,��׫��)�2,I+~���(K�*��'���5%N�r	����AN,���.��_9#�j�;�v�bh�xJq�ᆠ����L �z =�c��E�T"H�k@(Xrl��}���O��Y��Ā�4{ '".
t.Mu�#�ʋnkk�1A�ÍJ�s���YC"Q(�ԝA�ӡ<���X���d2f���	Q9�#P�����D��qȳ%GM�����Kx�Q����7WO5�C���$J��mx8+�����w��!y�o�T�n0��6<-r�Z���~y7�� T8$+K�6�+����93�N��T��Z+�:b��F��mϛί�x��5����|����ו��?ip�wg?wx��c+y��ƽ�W��z�t�]��O���
3��Yf����_n��*�b[)�����"�E�U�;�"�D��5�������ɴ}3�0�7�s�����k��]�	�X��Ώq;��7(|J�6F�"��y��dd;��#k�'p�n��M��w��+Y���)ځ���;�4j����#�].���/݄�$U	U��3�,z�vic8�E��_��*��A��&e�Y7) C�x����}�z���sٞ�����bblj�~��"�[��g���o�-��YYY�R�(��`�	��/_�(݉���5
o�cƜ
�v1V{8e����3�y��������ó�����
��%����O��-/��-��$bN��t�� 
�t��s��D]B�Ѝs2h	����U�>yBN��� ��Bq��)�t����"��qBC�hu�iu�Nn�'|�S��F��=>������l���
Z��HJJ�(Q���~��+��[�q���3���V`8ۄY�\�S���&���A��}�h%Z��l���'�>}�7�$�2�n��1�h+2��%N�4*]=?�������:���w�(U#gy0����sH/Ѳ�omC����	�.m�3n�պ{*.(��n"���=��Z�~@�1�peQ㳍��F�U��t��9�,9��SA
t�8ŗ��##i�I���aFg�F��L{�������Uj1�"��ǳK�=4]fs~�֯!v��P�F��6��;W(���v�Ͻ�jЄ�0��s���,%p¨7���>ʱ<ϰȬwaA�O_:��|��F������5�vJ��5e����]5�Ϗ���5���J������v�����m�N	�0����G��GiiU��iߔ�?�/S���Z����ro{�r���me(:����;�Z9���Ռ����蝜��;;�pG�GF�$f�҂v��<h���!������E��[������(«a/ �CB%��f� ����ac���Τ@�C���(Ƨ����� M�W-���_��^P�L��X�����Ӯ4�حO��9BEo���d���������?�X����A�BCò�ڡ�Kk�����}��l0�QD;E������x�L����־}���3/3�i5����m������!�
��+��SN��5.�gy�y��q���X���-�(����G:M�[�h�/�3h�#[�:
t"��Z5?��x2�Y���ꤢ�{���Kp�yu,nWd�B�8-��C�٪x�;�M��#	�.b���5r�%z����;�lyiiԟ$`jyǷ!F�9i��&yr@�t��g�R�N���Omй�b/�Ϡ�R��"�.,z-N���U�O8	�V �a�©^�
�>�ڍ��>(�V��%;�75@5g������!0�U~�61���8��u?�lw��.ޔ��`��h��di�
�63��1X/.6��{�� u���w/}�7�<���k�����S����*iG#���A��T�=y��јV�ڍ�>b_$f�@ّ�����h����C}>��^Y"Yf�wx�B��t���\�<@NwS7<jW���S�7�J�	b�%�k��p�IpÉvНsR:��3M͎)�]J�M?�h��\k��e6G�?C����a]$�k�US����M��4�ڗ�l�M5�h���V��N�T�]kx]�Q���4��*c
�g��|<c �k�����W�J�/���/o�T�u�(��Ү,���kV�St����k��f���Z��R���#ʳ��(v�?5�\�c�X|F��z���������݇��>�on�*<�"�Ku�[����I��7t��=�[lfgf�p����p&�Z�mOƲ��T��6��1�h,8�^>��	�Ң0�i��}MG�I������̨z�$A�`�U�(P}���y�q� uH����  c�IA��M��7w�ړ�1/�v�C'g;���F�7H8 Τ�I��Ih�����VaC���-u�l_��ٝٗ�W����
�|�ƮP�j����1Lx�Һ(|Л;�I�%��k����;���}�k�j��T�ڍ8��br ��4r4}SVm����XY�3���9�P���u��^���c�tU�Ӈ�]��b9�}��V���6��ڰ��07Zҿ��T��_#�p�����>4^.n����u�w�A�"\Uov�.��h���0��>������6���@3���F��b>�(���9����-�k1�Ԫ�R�fT�eI~.�C{}����3�+5C{7g�����@����o5���0c���KM�[	ƨn�M��!�~��5Ԕ�Mh�:�<��{�M�ܐ]��k\�¯�t���ѪhoN�"z?�w�N�����T&�/^�#j�WK��j� �a��-��nf����;Q�g�9z
��n�Ãs�K݋����l2Ko.���A��z�U�)ܿ���f���*�s�Cae��L��q�^�O		���y����:��D�����|~��L+��f���@A�y�����hj�N1ڗ�X;OiX��1!g�؏T-,\�i�|�2x�S��i�6����]�:a������?5���כ�� ��!��Z~(��U���,�X�`�@�.;�w�PrR��8�k�u����o�}�
�d�P�N��X�-���f^��%�7�r���Z�¹�����C'�$C%�n��+T�Y�n� :� a3��WU�H�A4��K@Ԩ֜x�Xd�B�d��C�⟩�������m���ac,9�����m¸���-*h��^A&Ī-��fͣ����J
�,
�5��{�Q�cZ����Z�:�Oz��q����}�
�������|�WF��;TGք��m�q���FI�KS�!G[l�R����ׅ,�tn�s�ʊ�Ļ��6���)mMM���ߍ��K�ؙ�4��眓=��V��md$�ǩt�QK��?�E��2]|)�������5)��q�t�p�C­��ԡ�
��s7Z�+lH.}۩�m䏿������30(4���r���:�. %G�ם��%]�{d ���h��^�`R�TKS�5�#�9p�7�T�ϸ�IJ��!�������?'aD�h^���}*���Q(��N�*W�O�Ҷў፻�Ka�����+4��
 �ne�CG��#����� C<\5�ۏY}D
$�Xsϰ���;���T'ϑ`9,�O�TܕP��8լ:���%�E��eg��}�ϪR��Se�7�;��UIb�kk7��&��ԉ�<��U�b��z;x���N�R�3���=���L4<��K�8ǟ� MA����c��|į���ҋ3%�@ �C"��(�
F��?��6_^Y��b]i�����ƫz���^���
��>�Ԋ#TT���W���\=բD�k1�����o���g'����s�H���N)F�Ȓ���:F
(�Ui�\��]%V59���
 
I��k�+hgG,�h��M���-j�Ū^�ؠ]$|�4��{�C�tzow7H��-������	`R�:Hױ�5Uy�	��	?���B�Z�o�5��K$�_oȱ12���eQ*F���L��`�~n������й��m%c��2�nC�1s9����:@T�����s?o�bB�������{�Z��=D��@�-sFÆ���J�Hm����]�Y>D7��Q�t��d�#]��My�E)��m{�݃���s��I�V�/��Z�0�E۪l�4��?�"zv�4Ԯ�L�ܺ)�a�p �<���F�w�Sn�n����e l�wN�vPP���J��źK���&T�8�gh��C��iW�NL=���h^On��O���-��~�Q���o���j#�DX.+g���o��ɗ0���2|i{���N �!����|h:/~=�C'�`U/�U�]7�7.d��Q_`�Vگ��E��/��|�n|m�9�	�n5�FR�Q���Jm ������-+�q�Xk�J�m�#� ~j����HdHش��b"@�
'��YT=9p�\2U������yhv
��і�YXԕ��_ �z�]}ȧ�W�f8B��f�?�� ��� Mjkk������Y��}y���7�î`* bX�h�Q�$u�n���Cu�!���V�!I|(���V���{����J�$�s�x���8z@|m]]�ΰ(�fC�%t�z��z��/�޼�]�� �\�\�,]�6\��Qw�gp�?j�d��9Eg�>��YMؗ7�.��%ݱX�\��XT�%��(�/`��(wfkk�40G�9B��?�C��2�X~�\���*Ԓ/��}�]��v�a��U.�mmvG�0c�ڙ�Â-��V�<H���6aw��G�ڝǗ��.�w*�%6[{�m��"?��Gfe)��.�R8�$gx?G���|;?%e8��PT�Y[/f$%��8��޿G��Kw�F3��|������E�����PM���O�t�2H�˯]s��#1���J��P}/`PWk$(�v�G浵������j�Hf�# <�fgmo� #=���M�����\u�查���3,TF������zJ'�fV�4	d��Ɔ��?G(t*�7�n�vt*��	D��/��+<�_�{qNyr����b�1��*�Q_�[�@ɝb�c�������P#D�^�d�404O� ĴI��*~�r,��t�*v��#!G'����
�=L��mI+��g-��K�c�� ��H8Vh������Pҕ�RC�LP��fP1�%?Z�kn�~���ՅS͊� #�X�ud�(k�����[�98�,ȅ]�% u¾���� e����v��: �&��JpK$����|W<3�h%ῒ�Lp��48X`�;����	�(���a��Ԥ���hլSmN����.�h�j�Tr!06F u���<��<	͋R�_��LL�:�g@Ӣ.�Hzx�^�v)7fأc����� 7�<����|�`|i� ��̴�Ք�@��������&���;����x\�i-T,��yؙd��=p�(�^2Y��u�U7___��U^��Uk�)pZ�#�fY�ޝ|����NF}tK�a�ן�i���-���d�P U���q��������kE��

��N�pg��o�7|��N��ƕ�L�bE����D"�ɓ=w����𹅅�x��e�6F��-�>\)b|�#�#k�Q�<GhT����t�Fj�b�'�-����w��Z�?P��Bh������;��&z���+�w�Z观**^��#;��/�ɱsm�7ط�hyi�ʛ����18����
d��1�Ċ]�����)�ij�AG�>n�h��!^����s!�i�U��������M&���G6 t����g+޲q�e �R��3�kg*N3�-����9�k��������_CB7 '&^ �6����@-��T9Bٔ�lV�{<��\*����HW�]����`�t���l_��iP�ڰ=��"%U`ꢌCV,o
��՚\/u�} ���I�`"*�$T�vl�B�D����Y��#�k�}���~2����6��1��w��֏�uww������#}��q�=�ov�����m�-Kcg}����J+9e�����r�L�bT���L�����;{��uw�����n����UV~�z�Ư�=�[l��8���X�x��M�M��=��mq���ӿjg� ��@L{�/(��#B����ʽ:E�z܅hc�ĝ>@e&&���~4ٵ��	�lw��F�־B�	���tgE:����p�h۬޵e�rc3e���v�`�j�����2�<:���>���9��d���#!��Jl��&�����t�������`�3������o9��iQ�	j9��1�'�1�����"z�y�4���_Q�����{ĳ�~#�jo}Kh:�3���2677�l�� P�֐H�����qS���?���ݟ�����&��QW�~B�;�{��P7-�mycr!��71OJ�0[�u��N+����֤����`}>��O�V+K ��ȱ:>^I	�jR��t�n��r�s>�ʍoL�e�zI�^�#�䤧���3�_Ct�?}d?�@�,~N��Yh.5�1�����o�� ��wyܻ[tyI���v�0�!��-*��e�(�}���|��б��k(6�B��p�!�5���s\�gz<��h\�lܰ�j}ܗ�t<��5�#?��XcSA�a.v�:ᐲ�������:�&�ݝ+܆���������כ'h�r�B��1����hAD�	�͢��)g"¾�@:;�{x�w�̚��4o������`o���lj�[����8���Y�]y���%)h6�m6�a&��z�f7n����Y��ڞ#�%^3F�5�.��뚘�M�VJ��|�N����x�<'g�e�
�ڸ0������heuϒ�z��3c@+A����lB1��b�e�Z]s�rNs�c�������:m1cI���+��;!I}񥓢�oc�?އV_�g���1�sQfg{�����k��J1��x�X�����cSZ|�İϕ�[ǭ
��́��c��+� �[��Eu�,~������T�<��C�H��@��I�vk%���G聃���'+&�f���oj
���]�4@a����i��Ax���˖j�j������LLLjV�A�����S<���|Vw��l�b�luzp���ѣ��g)�;��K&��S�n;f�)����Ɣ��WIM�2��c�N�K!eP'$@�6v��`獵���P������#t��C��n9��>8%/�Đ��P��e}(��y��cX��뾱��}�,��Mw�ւ�U�jkE������C5��V��ho@? ��ɩfc{r�bF�c������?�RA%zhӔw��Z�M2Pu�p\`)ewWd����S�X���P-��]w g� �zM��ɃL��UT��ͤ�ٚxchtP~�66F��&3ǘ�Vm'��X��la >���8s_���q��ͅ�����Z@.Z�(ѱ�����o��ola�[k��|JLT4�~h��-�ҫ�=T�B,�9�g"ى�e�&��2f;�L`Mdl�����L+�����ݟ��+*�RN�^ˀ��d�������ag���@��@ޑ���P�
�v������$�#��tFWo�wWP�@gy��*�vTy�C��.�c4<3���ʹ�vsҁ�^�xʉT1Ћ|�ľ�؟��#"�����[D�i������=�z�����g;���H�ӷ�|�b�����+��h���1�X�ʼ�Dq�]���Ȥ?μߧ��k�	�C��&����o�Vy󹊖���!%v�����[*�U�*�P;�a S��h�Ym���w2#�����<>����w�	����$m��?�i{���E�����t$8��%y��Ob��\ll�O	N�j�.[�ݲU1%���/h�s��'r�T'�����D�]��<�>k�'?�~���꺕���Onu�&*f��$���a�?�ح[ �%�� )/))X^����Y%J}�mT���:����g��/�`p�1����)�W!*���u��CY*�c��rZ??&���8B#GLj����83t�TKKIؗ�ݫ Y-l�PIJ���!�n�UYD��8������Ą����i�}��y���0�諮�v-�Y�c����{Z�Z� T�DG1�6��O��?$�^Ze�O��k�[
�$�+$1M!v
� .A���DW�C%P 	�pHV6hqߴҴ�B�u��Y��l�8zG'73&Ʀ���ZF?E�¨UlD�rMX�r��I>��n���.��㛾c_8��=幒��fy#���])�I���T�0$������5˞�ȍ.���Š:��>p�b	D@O���H7�>�t�N0��L߳����^���u�� �cwT��G�����e��m��e}%�ɲA����09�,��o(�di��C<�ַ�s�v��=�?=\n�~�z+�~����0�G������\��\" �'m��r��@l��^
z�7�3�}�< �=d���`�,&�Ͽ�ȁ�A�qB�g>i��?�9X�{����sGGO@�k�]:։����C���CK���c&b:^7��x��B�҃�>��*�j>�%��,��ω�zh=|��`|�CB�?ڢ��w[K<W}���+.�����͌3��������ҟ�7�-�'�I��>"�=Բ{<���Pg+�1�ogGDh�S\�)9,ջ�ig{�F�
�H�h�]v�U�FA���^�<�Ψ��A�wY�����Do�@�Q������=eD����T���\�n�bB�8�����3����#q_�"@VfeA7O�}�TW���5�_l7�aqj������錇���Bem���jKLk�{6&%-`�xxx�-)Ȟ5�Af��_տ�=Z�&�{t�k|�g�=�����R�^��MF�bu��vЀ�1���ɴ�D��q���Q��Ҏ��=K����67=�Zhs �.���s'}���KG�![u�>Q��]��-���G���$H�+)x�(���f�(��)���Rn�w�)�1$���k�I�մ+\��:�>}J=�u���;n����f�� �k ��x�e� }��h�N��A"�y � ���1lw��Yj��u8���hC ��O	�i�ӵQ��&'��o7��nL�% ��rs����n#ɪYPPD��A}��� �N�:�b헀s�4���3Jw(!A�սE�\��?`��x������nx��72};���w�I���c������x5�S��޾�F���E����t���
3`zQ�����o-I(��8`lf���P�2���	��q������i����C�Y8.���Wo����s��_�2�Z���3`�<��������n�ޅz-���}]]��� �{�i���F[�@?�R��7'4Z�)���?G���g��=�ˁ'v� IA'�?a�JV"�.��c��p;������H���L�c�ss���x�Ԉ�x(������!9Lp�;�ZRR���Ϝ����s�I��f�5���{���ai�xp�i�����WJ1!��������������%�<#���AA�v�m��"�.{ػ�j�=��BE�:F�]H�����?���0�P���[d���N~���M�[������U���A?�1�$?���^�X�&A:��(Vk��0E74��'ï��.*#�����;�U�n� �j��"I��9ձ����k0ļ�&�И������)�˿tsl8�����TyR2��q1��S��y3��9�������dp��=x�\������}���#07	xE�6#����$�r�S:{��j�����;�K���P�9�1c��Ǚw.a��ۿ%u�t�(U�>���Aii���+� �UBJJ�����߱Q4:H���?��@�����IHJ�����3}���&Tp����Pu�9���7-e��h��1�}Dp/��N��"%&Vh�*y�[����ڻמcM^bLi�,��_���α��{Ȱ�#��$ov��IIe���d{;fbr�������'ؒ�xQ7�;�
{m�#���4�՛�����6���Bܵ�H�r0��/���!��vIW^�v�� g@d���e�P���" �A�r����\a�f݁2��3�	�I_@�/�߽���(��wm�����F�	@�D�:B,׀�=x���s%�у��Y��탶�l-��mHf|������j�d/x}fH��:���4�������~^��&˽BB..�~���aB\di<�L
lZݢ�-g�lы�7z��I~�g[��o�y������-�
��@��w�X0��V�^5�%�	��j0�� ��2��{���������������HD�t�޸�,��������ő��ِ��f�9fL"s&��Z[������/C��<���~l�Q�-��,�=(r�_ �媭oI��_w�t��)\D�#''g򂤤d�nw�K�1QI	��!=ՠ��{{>��c�x<�[��[�
�KU�C����/��)�;K�1�
���A\��3�+��� 6+ PMW�{zvVz)��Q���E�:�!�O�� Yq��Q7Ru�	O�&%�h6'I�[^��bKٹjSzpe����IJ�٠��鐤�r���hxxc-�/(�y�lw��B�ԩ|8�A��4�����9{DD���x
ԟ��Q_C�1C���f��15��<���ql�Qٵ'��������������0?>:��۷�P�����[����#� _�:=K'����+��6F}�+a� ��ˍ�: 髞#I4�����]!l(�:p����-�ye;L�_�¦$��f*H9��|���Sa'���δZ�_�)���de�����2eM7��x�U����5�۞��?Ѡ�.V��RKl[�ْVv���,kf��8$����y��_Y��Qʱ"�7�/N�P	�����.��1x�g���i�F=�Z�� mѯ�nzZ�fym���=z8�|&���q9"�k@q��}2����e'����=k�1��ץ͔�o]j��M4燹�1q���������:F���,Zl�wh�����R-�n���F����~v�ш	�X,X���5�z�/B{�Ą��ޣ"����\��K���� �Ꚛ��$�`�([9�]C����RGd� `�}���A�}������a�`D��F��TG�V��4�~�����Q�d	/U4z�� ����vq�u�n_�O�X�a��0&�fA����
`%�
� �A��[;Q.AC*�Kr�ah�q7�"E��=�[K"�����o��ꈲ��z�9�f�O���Z�h�"���'��;xmct�������Fi��޼��T�\22��\�k���n�����D�2Xē��e���i���:�[��-����H��"�چ�Ln�bm>���Q��y>��@�10ЀJݯ����#p��GD�P�L��O_��u�Ի�p�v��F�T
�Yx�M.�/f%k��|����\?�/���pK	�p �-�V&��j7nY\=���\"�Zs
���٪���
����B�eJC�;��0�=:�L20(;�|T���u��l�\W������a�<t�.axd.Ĵӥ�^6�������Y����ڸM�3"� �P��f�Bp�*���\����S���:���	ך�{tp=qp0	�(tƫ�Z�ʼ2<ʺ>��d l� ���%�_QQ�U9/&��vy�Ѭĸ7��{<�T)_��ۗ��S�5e��t\��s�ӌ���oY��d�����?x�Ů�y��S���%�r�Ue��>��p��`�0%O�ɍN	ڎ}ӆ�|ߤč~k�)q���?�R�9C�]�z1����'�׫z�q�l!4������l_"=��3Ր]A]��d1�n|�YVkMsn����I`��:%�mX<��$�J�t�]W��4�U�EwllL�k:�T܋H�6��9V�&۝���)����R���Fkzxx��a ����$�#q��9���@N�1c;�Ph�	�b'�Z�m�w��j�|����d)_�ܞї������pO��8� EM�$��j֚w�4���T
{����W]���~ඪ�o��\�鮚�7�:|��P|i۟v"�KP����mn�WV�7�5䏋�=='�ڵ��L#	�O����f��'��I`�t�*z�N���xn`D��P�7Ѕ#�4����H W�����K�ʪ� {"�{��
�v6}��#�|�e���ۧ㳯v��M[݋�if�ǵ6���p�����8Wk3��<D�#�޶N�k����ШZ�Y�|��3
ڙ�#�,K_m�C�����j�ҁ��̼t���{8�lvV��6�E�K��N������o/��'|��*n�\���>JY兕���dV�H�ka�;R�Ŵr�Zzc;J�J�pb��k5����`�����0��`��)�@_^����EHp"�$�x�Ʀ��v��msɌPL��/���S�8�`-���:���=d��gR
"�;��9�w�������wqP��C L�6���]<���v��I�h<m�JXƾ:?wwU���(�yOqq����2��(L�š@OV��R����n\⻎�]~��OT�q�!U�{�bT�V�(�۩\��;�Ǚ�Ha�l+��)��պ�I9<��2��O�ƞ����UJE�#$e����\���cz��m���,6���~���]t�/Pbh�[���g_ZG̙���uȌϯVYme���*��������g���^��"�B�Ԗ�x\z)�o������c�w�9{۹����ʅ.%Ͷ���ZK�*�o�W5�����M�ޛ���i��Kwy�څ���7�MB���P�%�������6Ck�����a>P¼���_���s
�]hPk�#�=�I�a�d�}�`{I��;�?����o�����h�_���Cx��<Sh��{��<�|����ⳳ���
���t
[ZW���4_��Rv��mv�)�O�e60�2%4:3AUk-�E��e���:��@��كG��[K�	��.^,L��f�n��H>?�L�Uou���O+ZJJIH���R�]��l�g�[�D!�}�"KCI�ck01J�%�c	��6���}�.W\%s��>�����rP��\�]�F1�f1��1���{�*��Q�ϛ���o6@pfB��n��:֬t���9�NGEG�WkYL���kk뤥�
��
�)?�$]���9r�Jd>��FR��-=P\3���e�~zSh�+�h��d��).!Q�������:�yI�{Y�7��`�� ��,�� +|�����u&�!"\�����5�-���_{����q�:����b8�Q[���hx���;�(���F�H�1Xz��9��s�"�����Һ�.�
Hv�������y�����`��#�D�V0h�Z ,�>��5��(K����76A��@���i���b�X�aVȢ%�N����Iw1���t�`��ݫ�,;��̻�[e�IT�� d�F����b��qɍ�K�"���]ŕUU��-KMK<���1Yw�y��y���7+���^�!�t�u�
[#7+�����G[�Ui<�6G������^�5jVἡ� K�T����1-�Õy��0$���/�l�毰C���� �b��������V��W1|mg��^���L��:^��h�/�w���,�|ͯh�N'�Q�ւN�P���=:���q��Z:Y��o���x�g�,|9���]`�������-��
y�=��ME�u�H�m��|mb��������B�K~b+26I<K��4{�ۻO1�uX�J��Ǎz�+y ���$������А@�

�u�v�. ����Vy���.�Vw�?�:+v�������ՒS��8à�\48XW�u��ߟ��$t�z�}�~ e�߿��`�𻤜xc���^��V�k�_��?ج]:ӎ1_��w/��ݲ�^��w��
>?쫝��m�c����/������=d dT2�pG�C2��s7���˗/�I�G"|b�&��G
tX��v����3Ul=�����뽏��Y���G��**��hu˭v�����|�M=R�+ ����g���/ķ�³��HW	@��E����S=�<W=9h�������p����������I�h��1�e�m���F�U*���~:�� |N��^k��0��g���]�
�w��Ƙ��=��r��Aj+s���$�	�_���y?4��6�(��%��C���4��ۚ#�ൔ�7gR�s�V����c�/�2m���󹕿o�����%�����0��36�hE�-�[��`-2,.�oWc��x#�=?r�w�Yk���΍���q��9�.7{�5����h��B��]k�Aa�����*�ߚ�u���*��|�����R6���xB��$��g�B:l�[���%���B	�S	F�z�^6��b_�G6�ȯO[���)�3R�<�����2g �hDF��?T�=v��۹x����ju�T2x4���We�{狅N�Y���q�ji!vb5+N�%�Ea	�X���ג��
;���jp������.��CϢw����^h�k�)0(�	�����x��%K���>T�s<X{��&�sސI'�d��8�/��K�z��Y=��w�}r �$zJcg�I����i��q�y!���:����5��p&��~U�ǫ�˼PMk,��x� @8�z��iJ:�J�w^9z
���Y#�����"�\��y�����h3��Μ�R����|������ʷn�je��
 ���Z�L�d6��Ae�AL4�]rnkٵ@8��`@4ud;�%pU<��Z�p�X8s���Qd�!d>�]���T�P��
r�䨟[z+����~�7k���'ૼi!1��>ۯW7��.e��d���g���y
	���Y;x;��%\Y��&� ghx���v��X��Ǫ���qY��dt!���_�<�,p!W�)  �7v~o�z����c�*��b��= Y��4�ހ*�V�A�tP��3����T/$���(꛴�膺{)a̍���[��F|SC?�'@1<��ϱp-���J�a�'V�\��Yo���y|�Y�����J���i���'�̑� �rtu���I���2���o;Mn�eGG���X�{q��牕=��J-9�e����՟������b/�L�+M���Y 0�����v��7�h��?1�W�B� �ƒ94�}|���ﰘ�!s�3Fv�#�p�E��p�� Iv巏�=\W��3K!$�p
��+{�ĉ����9+��1#2��$[)~��W�졮�Wl�E1��37S�{��l|ۖn!Z���7k�s�S�A���>��{n���ɦ�����f���L��W�ڤ�\\\&��Ft������WQ��J�fZ�9�V0V��)�]��Z3��;}?�tZ~f=jr��f:�-�+�YT\����/�g�U+YWhVS������`;����|�s�}��lVx821�f�#�",��.�/�0^,��ƣ^����;1thb'�%Z+���z�0�;��\U�p�Ω�1�F�?K�{fsss,z*"��W�y���1X��l���g\--���F��xUF�F�cU�����!�?�hQ��R��|�t�!o��諀?�ƾ��bbb�l�0�� �2��ʗ����Ɵ��������(�fWś�#�ֳ�g�;5<%�}��P׈��I�d9����7��=�bo�>Q>�����V��ipAn0�IB���+�K�-�s�vv�]m(Y$�sK�����ҹ��/�S6�ee!�:�������7N�9N��R�����NRk'��S��Y���s>�~��N�WWRr���4nsjȊ� XՏL�țl�B�s�{j�o윥����d`}����G%�x�I��Dֶ�||�����u{"ӿ���,v3ڰ���}��5$��i���������)0�C1��h�^W=�S��s�O�c��>�H���gKi�?���4Zo��kk���e�j���1���lp.�����<�)��6�o��9L�+�B�	^�S���b{�e&����Q8��Y�ɩ��]���|�1^^r����ĉIj,[n������tڜ	��<8i��-&�m���YWW#�:�ܣ��*ccc'O�Y�m�`�I��&���Q�.Kos*�jG �D�Uz�z�����!�{d}v���Xl�7n[n�b��yT��Bl��j�͢򒷗�������]�3hZ�$��o��&�C��R>�=��FaBI���H����J�)�ɘ��>�1���APr�V2���?�k{!d�{��U�ܩ %�C�÷��0��QM'B����uM��1�Y�c㤵*@��ݕN���龆�r� 0^W�?�
[ܤ[��n��RFx�c9�>��r[�
�΋6tQq���9����߾��r�ȗy���	���o���UT�N�����'t+��!�@��f�n��j�2���iii���[0e��d�|�,G� �d�8$2rǛ��~�xc;B�y�!.+�]0N�D�_Ѵ�wRCN�v;aXPW�j�4�]�u�^�}M�/?�Y��<},� �������	�X������|xP|W*炏�:��]ڰ^!ZmX����q�b���Ą�F7ʌ%������
纉�t�C�V:mSĞc�Q��Dے�ox
r����~��/{�Y
`7_�|FBJ�w��=r�]ss��A3�����n��浢�h���wJ%ee��G�N7� ��t�����Ip���wt�]���C�b�r�0h����Β�� D"q�D��Q�t@*:��ܝ��)�~����"�`Y�|΄
��֚Nn�F\޿����T�R�a3R%*�u�oy���->��1~�\���!�P�L�V��k6�'oʰA�OO����N��t
��:�nIR�<0X����kǞ$���dوf�O+�Q���(����Q�\]��DS@m�\]���K�^���%�1ƈ��jv.]	$��D��ՄL�a�R]��ع9�T[��ϒ�)�d'2�{R\q���}Лڒ�f�B�X�����_�=����&:���6iE��@�K �[!`���0J�̱��is���u�q��N�V�$u�uvuu��W���}r:��۹2	�F���.1,F���M���B��@�2� �w&�Z��8�i��������?b�Ɉ�rD�� ��ԝ�v��2�2T��������U��z�L^Ǖ��޸$��舶�>YAV=ooC�����8[c�Z��C#�������+eD�=�5����!5@�N�[�5��V����qa����e��OG'�8{�$ H80`nʞ�YdwGn�w��XB��%)ʼ��%��z�-��Fn,��Lw����"�	[A�~�h�`���O�숱�*.���ؠ���=]
����sso�u�T��!�JK������F��z�P`P�W� ��)�/r�Gi��##C�R�.aH�0�����Z���%�C�
 O�F��@���3��c�>ux��� ��p����³��p]�g���Gk3B?ѵ!�I�^ �x����3T����f%R�L	�D�Ϸ�K_�>x���� �¥$5��աX��F�j�!װ�&u]]B���<3��ܜ���)|,m���$\4ʃsJ7-1���_�82�BE�DP6���"�(�47��B]0U�q�O\��B��n.P��7�.΁�4�n��͝��K&�X��r�.�b;��&5:�FB;���94��V���eP���4?Aۊ� pI֝���pq�����������2
�����ա��dj�ND��']ܶh��y�$�ͩ#Ҏf�܄N.�G,��y�ݛ�t#��E$��Wy��嗣�=�"�(�#}����7��&%����m���b���#W9��ss�E[�{C��8��:�	=a�w�a���,���x�ދC�G"[�k��a�Ļ];t��L՞��,��tG�Q�QMw���4Ҕ:�P�fgV�5`������ǆ�ZhW�R����B����9_������vuyA��ó@>�VihT���! �u򤽝�)`�?c7*��^���#��������Y�=�,�:<��Q���r�;�����#0��	br�*�fo��˲Ȱx�5-�A��3C�}���Xc��4��j$&!?����wᠭ+�Z�:$v�ā_��220�J��F��~ȓ�V�����k ,ȗ���,B�~;4<[������ �2:��bзA��9P5�ݘb���@"��{�QTC/'ǚ�ĉ�\�M`�pE�����;���T����GNO��ӂ�WMɫ=�Wq��!�U6���}��˔�m5�V�Vx�����?�
W�ʕ���f�1%�b��sôw���j~�����;�N-��Z�ۻ�F�_�^���|U]]>�� �7�'+�1����غ���D~qII'�bT�^���{ܧ0d3C�	Z�%V���{/�o�ٳ>D�H�r�T���,elV"��>��$a����Z(\OOOKK' ��~�r)��Β�fBN��*��R��XQ��h��Ro��+�+��\:tamm!`���i�^�w�} Q�\�և�}΀��A�^��i�.��g���b�v�R�by��Y4�%�lE0�X����G�d�;����m��%?����W̑R�)�*��"�oox�������䪪���Y�U1�=�T3�X��ý��o;�A�s 갇2�2��I̍��A�
De�>,�"f��U�B�f��S���j��0�6��B�R[�1�-.t,|�?eDW:�b����U��έ�Z�z��N2��^�����{@)��}D�e͚%��W�%x� ���Xu��U)���GJ�` t�h+�K�"�zNa�W�y�@�����7Q�̯F/ '�h�,K�w�6��ro�֚m��j9�eŭW�9ݽ�ָ��Z�����T)�f�b:Pd��;���� ��P��ңV�:�'��>�y_
��H;������y���AC"��9�K��b�s}w�$�E�v���� �@�&&%�n�Ei��Z�vގ��*8�����M�������U�[��r=��<]�U��̥�얒���W�6�:���_��텂h3+���k`���rt�QLZ	�<֢�
�[{1'=��֘��?��R'&B%$�ɜ���n�O!��f���`;!�%׳zBlP!^� .�?���O���bh�s0��l�Qa<ɓ�)X{�ռ6�B�97��}�h�伛*�b���f��=j߼z%��-�Y���r}}]LD�[�=�����5gMYv����,} Q<<,o+���)�D5�MTcIi)2e8*89�����k�&�׊���Agi�ʲW���] f��W���u�-����|�;i�?�ȵ����O���%G|�76�){�VlEӒ��Eʼ:c�j'�5\�r�1�G.�&���V'7k#>�������x��[|E�d(P�o|�����A_�B�����+T����)�	Wˍ�˧��������!<� �R�i%Q���#׽!��f�w�T5O����8��l�H���}����K��:8��|]�������*y�DG��CS0arrr�ﺌ��)N��J�,U{PB|H�mf�����&E��Ez���rF�ѥ�oĵو�cf�Sb��1a:��`N���u�;��;������P�:����fBۧ���O�f%Yn�{�޿��xd�������*$�Ψ�BO�����=���T."��
�׸���LG�{�t���*3P���$�`pV]��s�]���0�˗u�B;��d�]�\(�{�6K�6s���-���5�f���kY�b�,� �ey�l��uvVK�G��:� �¿|y긹j6I�{nr��nטo�\^^^v�{W{����X��W�X�K^ޅ�
��- -�u�~N��|1�BBB����-ԧ.?��v.�+/:::�\ZZj�"D��俗|�4�#��t��X�N��)>钘��V�&�=p��:,���1E�A��7��ʉ�$4���ri	ٮ�ЮJ'�N��PHZz��NMc���P�q�v�)^9G�������R��F^B��OL�߇�"3������Q!X��j��v�눡|#!����g����4�����?C����5���/-jX��0N$=��M�{�PǀZ5�spa��|F�ِ�Ƿ���?*<�m���Y[[���~3v����*םP|�W�2נ�?c�{9=����n�X괧�)0I��������}�=ϑX;���������`Z�'�e����"�Jl�!�����<�K�X�=R�_�����Õ��|�:]\��/2��Kt&N���GG��bp��zTĸjn3l�5�����b&�¢=||
h��1$�W15W׌R�WqcR�Y#���3�>�v�L�0��`�闒�1�Mg்	��C��T�{�W*��ߟ|�d�`�Dr��Y�̸��>0�$���Ao���4M�<m �<�F�Yx`��'� %D,�R�������1�#����I�j�ֲ�+#s��f�K <�~͞#�勼N�A��04���~���j���D	ZvcZ��w�eo~>��C�K�bV&�r;Z Y�@5�ֽ ��P�盠z���z��is�Z��(ă��p�f��� g{;;5�=����&�e^ai�˸�UDH���-1H�No����*^�Q�Xx�X���ɮ�}AV�(�ޗy�\{?d�v���/�$8���z��'�ڒ�9**j&W88�Dl&��#>�2�{���VfO|̀�jhiu,ME/}�62ʇa���M�n���;ς�	@_+��@pq炓�� [Q��]R�1�U�^�NNzV��Ι��O�	3(]�N��X
h܃�n�����S�vf'���ho(����\�S}Œ����Χ�+���W\����2o���B�\�C�����܎F>�g�"G�յ��=7s0�5fB ��P�u�l(��M�XmKK�Z�F���} ��b���`�Zѳ���5�� ��_��z�%w�oq��qٕF�&;�!lQ7���ַC�V������	���K�����[�����~�ˇ����x���0R�W�3_���,����Ӆ��\�+1�#�"D�����`>���LjC$�YZ�	˧l7����$&�F{~p�MNN���r�Xzt���j6R�m��9�����T��ٓ%d��' s�n!Z���b\иw�֙39ӂ
�&�� ������e0��iii�K�Z�Kssm�Ly�]H��R��xH��y{�'��b`���na๠:����7�� �#Wc���K��B=��G!�8g�@�\F���T'=j^?�!��)��Jm�qG���5^�Qb���֣8��ք���ۜ޴�n>�`�+4"�L	+�K4�F�i<m��??��8@x�'�j���U	ߑ-�HF]���4�9x�_7I<p��Zi��\=�&==��N���};J�	��ydE��G[��i/{=`�,�o�\�{`m�E�Z�(�W����a�z����3	30�6yb�?h����]\L̬5�8�˛J� �}���� P|y`:���k�u��!>�Q�uϞ�X��G'g���$��0�C(��/��m��zw0�^���j�|L*�8�d'���2�p���?���0�U��.s\Z�=;�;�<1;77ݕF,�o6HMS�)���t˽r��C��4!�xBG.�����bE`u�(2E`)������~�G��hL��q"*�%a6VT��T��o��ך�le�$�D6±���9� 5�.���ևz;.q�Ĕ�M^��9�V ?������&/: �+��^�cvj�iMM� M��|��և�ӡ'_D����A�03�ܡ��@��H$i���3|�����@����C���~�Y:Mc�ޱ߳-����s���?�N���߷q�!QL�`��ʌB��1H	�G����!`[� �}]"���:	Eɹ���c����J`���逬Yߠ��������������q�+�G��ب�Hp��-��.W7�Be�7H�l(Ž����3��ʣ��Y�w���D�p����=#��SW{��~Te9X+�R��>+�X鬚Z$�[�++b42=+&����NWV��&�C��@�>~��~�fj�J�����7�(쟦)�?~ �F��qq ���u�=xp>g��ۯȾ���p��F��Fv���$����ɞΔ��Y)��x����щ��ݺ�R�l��g��_=+�X�:5��tV��^��а��m��(�Y- D*֚�*]�
�dW��*�*��Y=��������C�?&�D��*���-�
2
|�~��F� ]gZݷ���W��pU������;{V�6���:]/�z{��;ϲ)l���^K�fG髨��Z6f����#�����2��$i�#���1�f�܇0'�}�&�r	i�r�Ç�`���Z��D�_,�h��̙3E��Z��Yb�p�lL(�R�Уߪ7�`)��r_E
[%O��;�

[\^������ʜ��/~
؁	�P�p������[�I����]�é�1�DE���yN�� �O�
��<��H��?^v�M��uŎ(�;F졘[��fFF5��u�P?��������� ���N������?��S�G�Bq4����h�����ު�����1��JWQl�-�SQɑ�j���LKg$Οp��#$!�TH(��w�<��IX���#hi�Hr���藯ױ��cRѥ��M�������g �ݚ�_�ܽT�D����!Ӧ}���[� j�9����e8����>Xɼa��K��)d���jg�#{i�Ct���҂R��z��uz��sz���9WR�!���لh��Л�B�[�8
r;2��p���ل,qfxr,(���M ������!uZ`��h�;�i��KuEB_�D^��{�0KT���@��؞㙚����ю
qq�\�I�%&&�?�*<�W]�W?�?'"Է�*`?=]0` лp<�ւ�u%%�i
%ɖ+xl�|��''����v��7z�3%�lT	e#��*�N��l ��ӎ8~����*�;{�ZX$5<�����L��~��tu�QfJ$-	++^ ���@�J������\���`��T||���oN��8�PPKM�)� �2��	�l�WV��P���,�B8͉ͥC6����e��Vqj(�!l�/>ڂ��Zrm�+�r��ґ�����ʎ�
뽇+ݶ���!H����<G���S���0%Ƿ��ب>X�sB��t`6�e�B&tx���XOONJ-;�X��)IdJ��z�b�����*f�y��}m�O���7��ACV\��d�	�:߱5b��8 [�?_�,�ޒ�{�����2W�R�ck��V�l �D9y���I���\���L�d?M�&`Ĺ��4���JA9z��F��%�`i1�rtv6����TW��)c�ӽ����}$�%�@�k��y ș�U��� ˻���-c� 7*j�\�;V���Ԫ�
�Ð�����_6H���R��8#�"&h���9w,���>�yP`g��7��X[[��k���w;���[Y)���H�C�He�\@Nb�i�43��:��?�s�AC$����e��f�e8��È��`�Eμu����iG�і(�T��u.�����i�fck�&��fi�5��	�
�#�D�dڰ�����Z�	�����y;y�!���D�ʤP!���'����}|�������q�ҥK̓n��6]Z�I�����������=:�_H۽*%�#�����?}�]���^�5f
����uj��&F_(	�i�]r��e�צ�kK��h����#�6M��ț B��iժ2,��������-h�G��/��Z��:�A^�piX'��v��������>��Uy
kN��� Zpt�Se�F���	��u��%mٿ���m.S�2\A��������;@Ę�p��^^՜/|�*�����K�	ي��D�q}/�+{N(>��1E��-�_4(6�l:���v]�(��72*� ښ���iZ#�]��xW�dM�l��D<�fX�9ڳ�=U�/��N��3��\�ٮ���h�?�*�^�.��>rH(i��pQ�Bp���'�PS���2v|�	cK�*@V�>~DP�$�?"�&'_V�때��"ǆ�땳d8�8��>G���������8��WKHHp��= z@*z�	�b���ǎ"Lu��5��Q����,��Aw~�Zy��x]`�}�����};�㡊��$nlЉIK{�G�fU�x����|�E:��?���͛7�	I2���3H###ˢ<Ժ ���q�DɎ��˧���Q`@�~�x�1B�8������FO�s�p�^���w"�NFZ��e>VU��l4S@6�����1?�J��?��L���?�Tw�A�ς'C��
�|������{`�Y:k$R�Ģ���GV�!VwwD�������C/Oc�_���C�T	���:���{i�mN�fG�H�l]�1'ln�j��N0rM��u6�����f��1�{G^M�xIG���>!�BK(��w��o��g�N�<�����	$xp!'�F�^"o$$"r
_�Y=�������'��)�XOr�����`'�H#3~���U7&��\Q��z�'��>���ϋ�b����Y����#YԲ��i��⋠�u�u����^��������VUW=y�Ϡ8A�r����9YYV�����+�"�8���C�������yS�!���愝�לi�*f�vU�܊@�b8R��+�Y-���2A�ڟ�Xj�F����zpW�RX�����E6h��l��=�nڊT-`��|o�e��ez�/0�[�%%%�9��L���t���*���2�V������y-�IG�ť}�N�c�O�F������/��>_�|
-�_��А	�2!�22��=�	��n�=�mݍ�5(JQdU�.#����I�r�{�#�9�Σ�x~��	��,@d�ǤD��zZAN�3����������G�1ފ�2d���-���v����5r�u����MP�E~�Oډ�?
����N�#�݆������]p+%�X�,/�������TS�=M���
@p۰�q�EAU�g��&7�M^^>K����2�����_�,P��K:*T{1���Ç���)))q����5�������?=�p������	Tf?Ƚ3�_2
���hAr�QW����#�����ص����X��������Q����F`}`�<j���-������&{�XCSɚO�cT熉�y�[M�h f���Kƫ�w�� +�2����f�%�s���R�Z����(��SEqT�3A/D-��H�M1Z����r�u}�G|�"{��%u���gFbg���Gw����M�h������i�Z�n�ö��SL�?���|rz_Z�Ҳ��)hx7�Wy�`��Ƙ��##�N..�k-��Y�����/<褔+��7H�@H����=���LD���|vO�^�w�wy`f��q	��F���]Ȇ	9�w��-�rv�8�w2��,��QO��n�h��oҼd�6=Pb:D$��f��9$��$aA&L ���z��c��"����S}��.8�*-��j�-��LLV�Pl�������ޠ���<F��	�T��:uL�!Ï����g�f���V��j��,�m�7e;�i�F�333Kϙ�95�!wq9?�G��C* L� ^L�2���\���nD޹o�0r����*�@���;�{�3�:�b>�e�����ʀQ�ʨ	�޷s�w��0��d}Di� A��<E/�!�E�!p)!ezj
)Yd��>�m����q"�+����������g���9��uy�eぶ���?@VB��sz�6��L�t˚���G�]���A�L�u^�eĳT�{y�Y�^�mz���R6$�9��?N��6�|7���R6eYn�gw�NZ������M��@I�2G=�����>̌q�Z`13J����}X��S�>��mYl�6�.���ċ%�� s�����{o~��R`X���CYn��TQd��A�](6u����.{�h>*cg�=�J�{j�o��)G3W׌�o�VnRZ9���Ӽqe"�}7Mپ3�q���'���=�L�J5����;qh��o�k�|��	�������P�+�puՂ��^���6���*1�Ť�#{�����+�O�W��o��iqW�=�L%�A�y�b$��b!dupQ��v��{gԺ�.7�E��{ڝ��H6v,�Tȗ`�[����n�A��h��]�١q�j��w�pOZ?�$��g��^�[tC��a���}���69�n�������tx�DƔ����9�f�^�2|3��j��[��Q�<V��>��G(�2}��<����¢׆e�� �׍���~\��m������&w�f:w��]��{+�o߿_��{ �]��%}����S������|�V��2k�^��S���d���r�V��O�S�E�*������^iۯn����.��X}ek��=p����~j˧āCD�P��N��~ԡ�P�&��t�gO'����D[�ۯ=�hٽ�����45�O#xJ�tĊĖI�Ǐ��t��u��a��s`�5���7[�y���W������Q��Z�XWZ��Ӿx���0�!K��x�����|<=�����&��)��Yk�%r��%�q�Se�7E_}���HP=���Fߗ
��ӷEm��V�������I�b�#�y�4�Cw���o/�X�4�R*i�ׁ�;��Y��H��ȧ$Yn�9R�5Y���^J���o��3g��5�DFvh��M����15�Z�?��|�c�m�� ���soǷQMee�>[}�MBr�f�&>^o��{[G�w����t��$����ނ'11qt�ǹ�v>�۷;���)��yxZ��T�[���{v�7��J��貀�鎃fBǋ��zS�<j3�l�}W��%z4�va��/��:�7��O^y��5LȚa��^�?��|���TOXx����p��p�7�inN���$w���|ģ���4��54��1)�~���ӡ����C�^�tH1o�r~G��i��<f�r���7Y�H��gEv�E�n_lcL�ZJ�����$�n{�|n;���ܼi��%vq�#{��~78OH���q{o�/�H<�5��td�����W��_3��~���}�Q��	3&�eY�5�~�$�8�|��	��k~���J〟9��m���UEDc����W���������?�T�-a&4s)V6�#�7t�5LgЬP���&-��f���֊=)�бG-�?�<��3���Y1(��n����m������e�
�p�r��s�'��=<8�3(&33��������K�z�||�C�,�q��س�|."�R3�O��9~���QX�Ya�'<M��Oc����g�,g�;��Jw�9gn);38x�V�M�p�����~����j�)��,C3�n��1�$�3#_'6Ϭ��&��֮y)O�N���@V�՟F��b� =�~� ;�^�cn�H�:C�6(`��������� �/�B��n��((:���RC�C�Bm�Z����b&�юU&%��sñ*Ԥd�Jen�#�ee�-,�k����>�����x��sٯ��{�2������y�u^>�d�f�
�:	-���"��E�
�b���E.nn���ZCG�������u,�����lN���BB�,�?"�I���Q$�:�WI��^�ɖ��s䟉|~���w���.�
��v�w�i�w»�ˑ�1��#�N�(g��uƈ�m��	HH�x�RK�ƨܼY��}
,#���o/������g�og���A��6��v�rMH���W�Ep>�*RY~\��>��CrRz�"�a������No�J0H�hCv�Ԩ)�yY٦�an���g�޽�����fY昹�Z*˰�Z��(&���y?�y�@�:��Z |��Q�&1��|RGA�~�p����Z����'��@.����P���N���@/��b���r+=s���@��������x��]�R��x0�{,e��V���9A�Ӏ���Gz�{-1�����*��V�JZ��������?�1�6(����x��ϥy�F���/� ���;��0�fBUR'�VEaG��,�}���I��w����E4���D�_�hI�La�ȜY�"��m���u36���ϐvXŧ��4��{�b��#7�;���?�7ND�k��hjI&W���-�ѽ��[���I��	�l��K���f2x��]�y�4��K����Z_bL]��=��1��dxee�8۵0lic/�\�1�!_�^�o&ًmmO�4�l.�!�q��:,#[�����ޞ��R��(���܏�.6�c ���n�U�LJ~����œ/�ki�ڞ���Fj��Z܊k�ԗ�xrS)�jRx�36�Ѹ鷵���nxj��U�54�v�%�/��Tn�Fe��ӗ�(��\���7��ך]/Կ�`1��u�X����w�o�~|��&�����k ��ॎO��О�yp]�qK	hT�O�ߓ�\��s�2���^X𙙥\�yb�B���ƈs���G�F��E���et[c�/K�=w���1Gr}�H��>�V�����S=�p��"����	��cimt٢̽,�U���B��k�L�������a{��������"x� �*�t^$m�y�9~2*��SCj� 	ʅ�~�
G1@"��uޭ���?''�!��mL������i�������q�4�������5x���z"d�A����q��C��Y��ߍ[�T	޾����޸Al�  ��!��n�̰T�j���HLy0p���˞���u ��eއ������r��8�x�C-d��H]t�a��fc�! �/V}3g��SH�y�c>9��2��ޛ5n��}w��7�
�jHV�w\|A=���s���>W��n@����3lwo�4"�n����}��Q<��ɓ���o[;;��k&���F�[�bk������W���~=�eK��6��Na���&pvu�����F���^Ʊ�����+Jm�}m���!T�qlᮣ#G��MF����Ǻ�}?m��t^�_�A��!���Ioh�8p8Vz�ܛ^_�x�78�����h7��$�'��?A���P��>�<���-��we�%�bv�"��
�������~�i�6�z�잣�A/Gᤎ;ƾ��t��%_m��+��,��|7,w���F�ł��r�ذf������ě���1%8�SJ���]��--��#��0�)+;��y fP��tP%��oa�g����ҊG��4X�n�ڻ�����.��T��Afp���U&���W�PT�7�t*���fW�f�W��ܛgW���@8������	�,m�E�苇;ǟ?� �me̪��𫍛���I"�ˡC�����6MO\\Kmn{��������ya&%��:"{�����|��B�>	_��;0�t��Y^���L)�T&~ϣ:z���D�\��3.7,�g;~�}���mR���Ǘ��h�f74�)����o���N��P~��nΡMsҿ��b��{�,J�&c�ڄ9H�#�8��0�2#Y�?�?����y?|H��ᘻ�m-�Z�@;�IӔy����;n�ftE���4��ue���q�{�oѤ�r�\ �K��Y��@�f�P�26O޿�x��|'�	OП�]]�2\O���z\���{�贸v���H�!��u�H:��y���+@u�	_��>P�9e�O��s����/���	V�3Au���+��|D����j�<��,�O���fЭ��)���ƬE�06ߕ�t�2ɷ>Jr����v$y[J,M���.r��k��A�ϟ����ʮJ�D�k��T�P�+�Q�c����>H�U��~�@o{�FG��eT�����3/y��t�3��u>}�.�s!�����.g��۷�G��0+>ZvG�����4�����xr�Pv�p�~P �Y�o!V��q��9~e�¢C�l.5d�=���U�l��⚬j.��'�;�т٦��5 ć�K�|�y���_(1�8z��;g3�s���(�G{y����(3,V���l�&��\q�~)��6�-*�� �<ls6*M���xƳ9���z*��:��K�ΰ3Y,���_�fH��py�}����>�<��	W]�������:��F�֎0���#�i��}�^erc�f�V���m�Ko'ڮ���؂#�y�H2p��z���^9�y4�x�ax���W�%u��R�}4;{闇1]\����33�ۍ�Y�[�ۭӷn*�?�~yY�*�2zW��"Χ:�A����$Z�n�h�wc�_���y���$nA�0��ks�;�NI �C�ɦ��޽{��A� ������S I�ըy�ϻ"���d�����v����y0�$���_M|]�E	,t�n�?�afBa�t�dOT���c�c�9�t"Z:jvVW���:�2%���a��1��n���X4��9�-��i�j���;l��QTt�e��\�X�h����q1���;O�w��"4��z���!w���4��Ю3gΰ�4���b%@����h{�@�&�8�}��,9t��aө{�7����z.�eq
?�y�e���x�����h$"�5D�	���D�����cbN(�����V��!�	c/x�Tx/$�������S�XE3!BʲߦZ�":��C<�c�<�u���>���2�yi�*ZV{��F����ҡj�����)��s Mi'/Yݿ��Q�O�!�W��jI��4[!�׭�?�������W	edeoB:���HBfFd�ʖ�Yd��|#�!��:I�W���������o���ܼ���z>�������z���a�%�B >�۲����P�s� �,� !<���6�].H�/�a-���D?&���t�$'#�@��X;8���+�������������թgOk���LM��ξV��ә�t*�����ވ�~w4XY����f0�S&o�C=;WV�|�����n݂b����fnn��^�3;3��Һdh3h��8hd�U��z ��0@Ɖ��`���++Hk�]�mo�m�(��B��R�o�v�ѣ9���=�B���qh������S�z�iJ.g���}� U�J?ԣo����tV343���~L%�thH_�����f���Q����C�#uѱu�;�`0~EV���{'��~[�2ַߤi
�/�֌Y:sPZA�Ze�4���x
 8}�+�G��_Q�uw�8nke�=����/w5+���X�u�ӕ5��9V����rJ�
d��_'�re�KH���$����f� 7�bx[0�o��X�m��=_��܇Ů��o�w�z{*��X�D@u����#诤:�ܔ	z��a�NK9@R��}V�"��M"��K��'�P�_q��J��&�x)$-��U��+3W���'q�j���9��a�3�]� '����g�ɕޙq��r�{�j`c�M��Ж�`�G�NWrWj�#�i��\*!!��@s6���==�GF�o�U�&]]��L_���G�3��@%�0��Ě��b�,p���i��{�Er�l��E�R��II?�[zWS��e@�4�(6��I�8R��$�?�Er��ru(W	2������Z�}Qq�`���Q���!��7(�P�*�ŴM���ݮև�z�G�1��Ύ?	�.G��!�1�_�O,��଴>Fs�H�� �C%���ɱ��)���2��,��� ?>X���a����;��������i�N�8@��v-+s����]�����5��ۍ�Vo������~Ŝ�Jӗ/ܴ�r�q]*��˼���""�k���P����n�EtN�⡖�`��}����R���?� Ӡs�)R^�>9��C?�Һ'D"1������m�MNe^�&�A�!�����ӓH:�x����Պ�ʮG�4jQ�3M�^��+�6L\�Z��w��A�k������� ��c��}�r>>[?�ǂx�n�ä{ֺģآ���@(�l3(���1�� M�M�|������Z9+�T���1?���[l�j�Uhϡ�L�Y�h.�<��{�I��'NU(�Nr���X;���%%E0YР'����J�/Ts����Q��5���8G�I����B!���({�ʡ���%��ALq�5rC�a��T�5�&�0��A����G��"�o���ᰥ(�k�1o��GoK<�L�Fw�8�n���\�%"ϵ��ԩ����mw߁e��l�!�0�z��ήT��gB&:3D>>����oz	&�g��BCgr�\'	n�TgQUE�֧��2F5���CN�葶7��&�̖WP@���P�d%+��Dx
���z�����R�;��{��ȯ��Fړ��АL��̮G{��z/

�n����om�����C�� ��͍��d)�Q ����r���lePP T��fQ�<�v���)����n�L��p���c��&�W:	a��n�6(w���"���U�ԭ��ͼNL��Z�=����k��
�+5=;��&姅��_z�D��Fcc���,����3���47W��]��NQ���i�&���KL>��i�9��o�iOOv8ԞԠ�/x��Ƃ�`�1�c��j�i�ő�w�~`�@��Q�N[��}��z�8�v֓=Q�����
�EA�'�pm�$edex���f��H,A�Z�ܸ���s ʟ�ΐ�N��#�:�n���}�'�����JJ��[����5m}���i~���~SSww�۷��~C~�SɕX'=`�Q��ï��U{�������>�뇠�d�����re�ژ�$�&4T�2���oj:ALӥ�<����c��!i�Ew�z�%��g3��Amm׵�[�Œ�x�d�5r^ۀ_J�K	9����=���R{'�������5n�<G����+s�Lu_9��wx*�
wG^^^XT�d�;���C߀:��E��u����.��#-��3�c5x�=��}9!a����
��ָL`j�M��<%�ׯ_��tjA0�uo_nϪ��Zh���f�#�񀋋�u=�x�wM*��%z3�ޏ ,S���߬Ӭ��*�KIO/(��C�,�p�P�y⌜Q�VO��M+�vVQ��_W�}�4z=""⿁hC�@)111�B��k�!G��9���.*ڀ�	���*� U��Qg<��F�j��o���n���X�w������Q����!A�0�߿�(�[�z�=O\�p�m�!M3J�S�� P�%_F��[/gJ����r��w��hv�}xH޽�L�!����78����cܜ����K���!%
x��u@߼��Ȫ�bpp�I��c7�i[��";��J�J��p�~�qe�s���t0�]����hy�,E*��_2���'Cg�������#u�����;��Z��3�N�H���٥�9��6�$�I�2Pdsϑ�RB�QE�R�7�����b��Ĵ[���L�l׀�ba�x���u���Z����,F�\�|5w�E��ő �_0k '�%��I@nu��� H����SS�2�%��[�Y8�|J������n��q��j$~�n�/�w���j?u�1��NZ���(o�U
���ׯۜ�;j��N%''�ӑR��#<�0��f��#;f�뛍h�M��ؔnUt�lgn��,��f�?޶��j_<%�D~�>8O�[����iJ�~/Ýә�������[�3��g��3@�v���'�|�B6��hÖ)'�����������b�٠HǝN��yҟ�����,��w��x��2;ղ�{Ɩ�Tz�����/��i_����ĉ<t�UKo,�`��h0���?Y�N�0i���6p�@�M޸��BT�����뢂�<ؽ�V@,�IE���V�j9B2rrS''����+��**�>�Ds`/��'B��&b�Iy��H�
����Éd|8��$O�(�����w�.P�CQ	ķo�Z�L�K?ϯ�<�'��^��Q317gM���Qm��6��JΚC�����~h�(��H�W2�x�@�� ݫ��� '��ۤ�	�A(�$'�t��֟����9�R�x^���6H�?�00��0�!�(��?�{{�.���UU'?On�Y�Y��蘵
�ڊ1���.:��gUqG�-OQ0q��g~��C{���kQƣ�R��(v�e��*�K�Ǐ�.ɼ����)���#��e)
9v�u�I��EJL���6+�>#g��#""J��PZp�<w�*\��ל�����erP�r1ErQ�J:Y��X!饜�*��>9�UQ��M�=<�Z�̫���� ^4�D�u�e)���gdp�'�L�L�"E��f�~Sܺ|�������*�?�
'��xv�d��|ae���0�\+�Q��<�/��E{\/c,�F�WԔ�7$�E��a�I���@|k��qs0��D=������{�	"��w��l.�KSQ��Cm���K��b�v)�5\��{b��z��靝WIw���=z�?8�X~�Z�8��@��"�'/'W� g�٨H?Aֿj�o�OT6a�Pd��-�/��䱛"Lv�ަ�������]C�FC2���P�f��*R���K<r�q�7������.�m�[W ���P�O�^��>>�,Y�f�����g�I����~f��I#D�A���8\^�t��Om��`�D�Ɔ�-w~�Bssw!aa��"�o��8��%R�BB���N���G��F5�k���Y�5�=��JJ�<~e!��
p��j�a��	�Y���_�6⏸T�^DTk�0������4��/#)��cU��E����122���ʽ������Ķ���Pu�d>$�������0c�3-�P4�3A�J��䖷�׎�����^��T"۔Z�l�RR���V��yc��o���_K�K3PQ*Q�I��g�4v��u��^ryj��uF�٫=�L���F%��ؚĳ�'�#�ﮪy\\&�����Vc������o��_�������s_BZ�etTP�bָ��� Ț�M	��q��!3�)i��\y�O���d�L�\��z�ӂ@i��ݫiBr���2�&�Zװ��jkq�81 _�B��5C�㿝�#,��x�7�H�`�T���?O�ò�(�>���ϺT�4B�HE�i+Mt}�a��tI��IIo�ּ
��-=�~9��_O����`�f���z�n�߇�BC�6%���s&wL���k�NhV	s�Bx��Urr0���ZZ���6ށ1jn���&�r�8�/��{��{_?sTo�����<���#��
׳&"�Y�YyA�s���R�K���~o���h���|-	z�]T���9�>jjj�jjN4	!R�˓U_�*HBx�b�[����'��2�i��pӅ�dM8��a��;����ij	�'7�F+=�43���&����dEN�=�_���b��T R�H�g��xm�}s��=#W���P6�Mn��p�ۖɕ����Zڈ�/
C�8��y��𡰄�EA�Q�DWV��ŬF&?���͝�RX �<<|C�5��g��3(K]c2߻�+��ݎ��l��v��ݔbk�����Sl��{��鿺J(.|�o~���ޞ�-:7�1�b@K��󒷽��t<�N�j��?/,�H����i�g���q����pV0h��j��H{s��Y���uI��⫢/�ZO�C�_�D��mF<�op֞��PH�� �u�GR,@���Y_-/��,U������8!�}**�i�7���w��d�Z�����������3��753�y?�M\��c���n��}�Qׯ#�l�� ���e�G�O��/ܚ��m�iz�\K �[*x}l}q��D��5"Г�����xx`u��F�c���f�Agu9J0�f��h(��ޤD�0E����P�eQ�w�����l��oo�����0���R�mW��kN՟��%
i;)�%�쯎�#ћj��^U��#橋o ��qI������.���iC�az�����U����[���tD	9FfQ܍��j}0
{�հ�O/;�84v��adѭy�Ԑ~�,V���f��ǠN��&6}�b�@��ɤ�-|�Z��`O5x[𧪻�E`L~��FDF�����5�.O��E	b	��� A�� )�����ڜ��~��J0�ˋ�����*28<�z�3z}]��Z48V�2֒�ΝM*2"�^��i]cc�kT�G;��K���_{�Z��N��Z树^Xڷ�G>�E��R]�)k��?�U>T%�_u|$S@sae�6_���f�ձ���;��G�ѥ���BBB$zuk�CdM7 �p8M���pӀ!8Az�"at+�t�A#;;�X@'M�����5&?��Űuc��Y�<a����maL�PJ�Sa����s�r�k��'�ĎTz�'�?�<N�+VZD$��n���r����1/��dj�<sڐ��l��a��iM%w
*���a�݆�&���[�!I�8X(L-,���$����o>2�04\�ܶ���-cX��)��?��H"��o�{my�~��izU�|���k׆Xx��	e?����؋o2�.}�	TxӉ��A��0�$)�@���h�e횅�����D�"liD��hO�����3~�彈bS��߹s�$xA�2=5�MJQ�>��Ī�&C�B���W�
k�Y���ۭ�n�չ�b�}@���~1d��?����BO�}b"&���yo�,mTT��iWrZaa�И����g�f�^�l�E
;+��@:N���5��H�S�P�oݯ��#����c�t���+���,���<D���U�^nؔ|�w[1�yv����빹|@�Ǔ��� ]�p*n�:�UG-,����_{��Ɨ�.\�1G��'��g0ۓv~�74;�/��]�{�$�)�LE߫���ZC���"�#9H��7��W˻i {�d�7�5�v�w�d}�@��L�T�O��$%%��'��<h�?��-�~$��X3&�'��-����& :_k�訓�Y׸y��_�J�͕Z#w~Ʈ^BY��vui@i�X��c�t����Z�)R~R�}~p��X��P>==�@%����6L�̃��⡶�fU��S��0���h'wN/o	'C=T�}�ܔaÍi�Y�#���w�Vn[<���/���˽����V������!��6qq̏�������1�OU���Pf� <���]OIy�)�>V��k���11T(��ё\���G������m�g�n&�R'Xfh	�\[�E�Ʋa~�&m���f,a gDDD���:�@�B�1>9V�{R�������\��i��6����Z�),��9r0�&$��	͚ ��KQ��}���������,$��"�z�֙���NwD	N�qE0.*�b%��0ٚ=!�4�ޟ��qt���!���Ujj 
[�b2����7���}�#�ݜ��f�++�
�z���א-~J9��GdYY�IRmӫRR7$S���C��>����N�`����j�iT�NIi��yU8hVr;��f_�H�!���[g�R�S�QeJ�w�CP�r���v֋�n�K�
W�>�m�c]�4��iҞ�\�'�^��_����7 �f�|�=_��c2&^��-���TUUA�L��Ry����op<�j���ڜ�2E��� ru������m;;����0��#�h�	J�*�)j�i��J}�G����7�-e+��;�}��suk;�]}���� &�a��Y�-�� ������C��]5$6L�l3+�� �Δ��T/!`6�7�)pq~># D��f�]���
ٱ�##`�`T~�@[,�VLݳ"`��� ݛVy�0�ys(A(,"��%��E�Z�h��T�B�Fy�X48J�Vő�\����M1l�{1��wE�2ńU�4^��XI�9
?՟��J͹i��r��/]��&u�{����J���A��ƺ�[�0�:�i��� ���L��o⽺ T�**����L.g&����8�7�35o���
���ne��0�'G��/H��)EZ�����1�(̤��*��Bd'���%d�$@���Y���1� �[�}�E:&��hB�L~e\�8��pexE�LBa���!�0P�Q���Fk�fO��~�C��sΝ��5��?[x�}a�""�)a��@x_�����p>��)Wד�D2&��'aP�`e���r��Rr�����Prۃ+BdYr���3����ԡW��U$x�7o3�=|L k:�*��EV�0��h�У��}3��,l�į���N�?����[��"��'�:{N.�$K�0v5��@���8͇��N����^kvC����Ca^��Ҍ���%�%�7�||�ݥ=[\�����+n�������8A"p����)(Î)'S2pM/��K�7eh	�ZH���:£�2>΁`��ǝ��Ut�HG6���r����ֲ��A�"˃tt�Bt�R������V�H>×ܞ2��rRc�[^��־��7��S<�fL���a��g�O�/��v7\^ZV���R�7��J�7L,��hl1�&���,ٯ���DȡB�%7�Bj�}�Kd]���u⑾84ױ����O`�a�˻'*�f��
�y���lk������3/��Iyo1�H�QR]���$t�8�Gcd���I ���r����9�7$3��w����Xv��S�`����;*�3���w(��p��"���o"��2d@��5z!����8o��n�D��@����i�26��w�g����yWU��V�'���%��`�N�Ğ�3ɓ����E�,��ڟ��|��L){��{�%� H��f�s�-c�n��=��t�����5���k�VY�`��C9^KM�3sq�%�U�־L6٤��V�Z\��̴�u���޹g�z�n=/�?���1�긿9*�օ��:.��1	a���p)
���TW�E�b,�9xӒ��༏�ET�G1��>7X���-���0�����ݖ�8s|���Q�)�`�(���-�|�mz�EYXY�p?����A50P����\���N�#ǲ����說�������]�!'kzt�2W��9����;���ڜȈ����BQ��['N������Ρ(����&�'���$k@� :��rP��Ʀ@!���s�I�JP�i~}�H3_D�ךۯ6�P���SE��J&X�[L��z~U,�)`	Tb����&�L�̀	m3�,ņв]jņA�Q����f���<fܯ4��V�Ūh��*'L��TL�k>7[���ih�w2E���j�$��6Y�	�7v,���p�{�����_uuQZaM�k�!��SNFq
<�w�=G,z��B���7ksČ������rmꇐ����Z��?	b��% �Pd=es�G�K����������H�U6�R��,\s5�
�Mlө��/S��/��lū,��a(���TK�*�Qة�*S��]��)xWR���6O���>8���J_���fY�Nv��f�cӬ*��M�s�K��iO���щ��x��0G+K	��@�j[ �.�U����ﶴ.�����ih#q��O��"���ϻ����s{�G�w��B��1�9����O9��%������>��Bl��8�M�[�������f�?�wo�Bp��_n�>�fh�.�kH��KD+(���W�sNUM�|7h� �8Y���*�U���R��WB<�m$Y���q�������?9��ҲxC���8�@���j�ӑ��A"?�1%���9NEjo�x�2��a$�7";��mٲ.$b�XH+ҹ��3aq���H�sT�iݓ�D���h����l	p�m�,����^QY������8�T�+�2T���������� �[�8#�<�g}B��#�h�����
�����}]�����Z����+Sɩ{� F&'i�v�]R��?�U���������Г�� ΰ�:Q�|��gqq�,ll�B]���О�ɬ�����Y��{6m�KNNn���7;H���ӈsa�"�X�X�8[W��\%�QV�$�x�c�r� ͅ<��U�k��'�D�6�o����!��s������A�<�Pup�(.ʹ��L���P��͏SDP�Z��К�}�I�#�O�s��_�z�O�|��e�e�VI$�{}�.�<�2�I�p<����{ך[
K	��W��`���L�������(eS���qZW?Q�GZ��%0d�F_W|��/ ���J���/��fWa.��뾱r�kt���ĺ'�R�S�|�VW�P�c�e?��7+��IY���,�LJ.����PE��!�~`P˽�������P���n^E>��bᑑ�R>����ݍϑ�'k�!��4;+�U3�/�	,;1aJp�y$?p٩��+��gv.:���� |1;�i�y(O�I���#������|-�XH/6�H����(�y���|^y��J���ᚡ�����N��Յ/.��A$�#��W�)	�vtI�yC� W�f�jО\]'	n��{�=���[����p��ӭ#5�Tћ��ڨ78F)��f���w�&�(2��4�^sO�ܟq�w�`��i���5�Gv�H��4��TWW��(˧�໕�*�iB����>Mf	��F��o�dJ��9����;Z��/��d��Xk�6#��/,�K��!���w�1E��fQ�dA#&�#Z)�����ץ�Ɇ�NJ�~�8�4����\L�{�����4 <2�;��F	�p����җ���qy�G�|\U5J��ob��h��%
��d``xn�ğx��M��9@!�Ӟ�W񺁠8q����@MY���kj��~��{|���aw�͊�Kv�s���2�/��P~5y�:����2�'�8n<�#|E��#�����󏍇��T�a]+#օ��\��[�z��K�ꍳ�ڤ[��f�ÌoX��;���$�U�?�9��V��yu�G��}��u(r�R���{>�2�ݿS#���=��4)g�3�̦�a�=%�������[R�o_��okm�t�D@������ͦ�4�k��榦��2u1�*4���%����_��2�4�����~{$��B�;?(D#��i]��\L��������㓧c
~Q�x�U����"��nP���9;*�~�Q��N��!�����V��ˤ,�։���Ndiha�/��~�Q.��G�X_{��Rbv��"�뗘�7e�>s4&'�� 5	��%>74�"c��n��y��K<n�]^�k����\�еk��X��V��%p�H�Pu���s�L��ڻ\�W��6S��+F��MSH#����e�j.%Y���%R��dr/��_����
��Q[W]�˳��YH�6!���$,	���-Rl&?�g�wԁ:�WGQ32Z�{����w�[����ǀ_�Uv�33��d�ls�j�
_��_)�b��.)�K��]؞ק��9Ԩ�1y����f3]}}d�LD��S�֛���;9�+e��\}�"��tpp���'Z�t<��`w�#�tz����|�bz�h�v��A��%8���c0�]	)�r6�u�`hy���T�A��pJ�� �|ᙯ�Ț\����aIXq����	�↛;~�ylс�^�ecg7uw�mͣ��
<yG���5�h3Ҡ�S.��&&&�01���a�N]�����J�{��=�B�0.���U���-?����meo��%6�7'+Y�Vn��Z�Ą~B�y�Ӻ���ǯcbR*�~zzv�D�T������|����  ({~'8�W"U�{��q �BX/ �)ϭwȮD���(���7jjj%ee#;�=n@�X�渋Qu�r�HI�!��W��ʨq��X��gώ)t�
Z��F�W&��^�t����V���� �S�Xs���%�*p�n�%Oת�Ɖ�(�j&R��0o00/:h�k���;�o+�!�V]�ٌ��,��=$Ğ'���E޴��P����+�����3U�;�L����)���4��PUV�ΙB����&��G6ҽ�
���F�bH�F����W�������D��_������Y&�=�-�@D�YkU�F����c-ܡ���x0��r��b;��#��}Vw<�(�`� ٶR�J�X��������Urr�k^~��i�)v�H�<k�Dl��O{jM���U#�~�:U�������m�����d����w���,�?�"�(��+6碨
:�!���~s��b�����I�����Y\k�����Β��RR�����Ƴq�+����^2f+-��{�URۃ+W��9eՀ���#�h�V"�B�ND���IY��;=�	GB�����aqQ�f����E�~ݳ��J���R]Bc�d��\(��~`�Zf�L[��N����^`���ž�a�\�+[�ω&c����@ϟ?/��跢���p�U�V�d���2W��m�Bs=��.���2�(�z50?�<�桴1o\KK���G	t��S�1�+f���z��-�����C�%##^�d�ݒ����� d�ܮ��L�H������X!��)��:��i��{UZ940z��KetO��pŀm�\u]��6n�Qo��Y�����'V�;P��[+.h��\�eVƖ�5��$X��:9��9��o��wٲ0�T�Q���*b������ܯ����N����IG@.�����<0�̭Bdo@x�sʾ�fB�][����L�X��t���>�6I�Ut+�����5U�!���~��[�`�_|��AKE�r�� Pm�U�᭣
�G����o��ZÔ����OB+�J����M"Yt�l��%w�T�A$������LD�f���A�)��gl��)�*<������RʕLL^�?5�	��t�MRjj$���(�P������N�:��201�7M���4]�e�K�Zj�� �R��tc�->��<S��LyK���I����,H]���"�U���v��N��T�Q���4u8��N(���5���y㽟�Bn���d�x�����M���y�����6�>�~��`E�������ӌp�	�������>�:M���_���i\Z�b`O�9]ӽ��3�~�A�9R��W<}>x��Lक़�4�݀`��>2G��h�JY��i<><�`Y/>{��ԓ�I:6�=�0�����G:Y{&��9�|ؿ��A�wK�L�����{7��zV�uN����K�ld��7�9kw����#p��!�4���ء�%OO��GN�/Zq�j����a�1�B������z�� =������{_C�����4�>�2�����AI�Y\|�ך����+��W�[���O�[0^V�98R��52e��m�ኩ���`0�!�u��,�����Y%Ţ��dM[�G�k�G������F���s�t�{�&!�J�g~�FBJ
o�/kЖ|�`aUj�ˍ��������p�����^��?�֢�˹;������@a��w�o���0��K�d�t��G��D%J#_*¼Xҁ��e�Z��*wzg���sK�Z�+:KC����:}���c��C��8�h��|-j`;Wz�R���])$$'�2���LS\�ڭ��ëN�J�WY��3IC���+�{o��Vfse&ɉ2ٸ�G� s?檃��s�i%���)�>��:����/�{k�$99YHE�Q�0<����|09{�R6���9��s|#�-�t���DT�����Y�X2��mB8E� ^PL��?#x�rq�2X����c��*�O�Zy�۫1�$�����ln�9=?���2KG���%��I�G-E1�����m�� �X����t��Nw��T�kkٿ4	�����
���`̬f��|�=q"H��%
$@�-4Kُ�9g;�wt f��S���2m��[:@���7E�a�3�;����&W~�.Z��ҋ�x������ Y���_� ��>5#I_���o ��x�9
�_&�/���mtO�2�L �	*w��U5jT�%؋�J�b)��(s�8}=���}M͵���Y$:KWVN����^Q�A^��g� �0�(��7�`"/'ssW>O���e������B��Z^�>�|���,3ٛ�Ib�++`q�.E�	����v�<���9Y���E��9'@G
7Mؘ@�	�	���}�;/�@5�����>��չ��L�֔�\0<�"NB^�PMqT.�����o�[B���U22;��Vp龍v�B=�.�;N��,,T�l6]H���\�,���%w�������9}�4�;$��K_�&q�x�D9VRQfuM���[0�Ohl��+�11���
G9޸����JJ���/䢻�9]��$�y�(CK���~�.�P�?-F~u
�;5U-1ND[N�1�Ի���15�_B*�$E��A�W9Of}+�[�LML��x�IoGEG#ۊIy���ee�	֛n�]�J�#l>x�#l�2����e�����j�N5#�b�}�P 1`����D�
�<Ea)	���d)�
�$/9¸x=��n�?v��[q6��jlu����
Nzu��-������&I-~W2��[��((Ƹ3u���J30א�U��>wf�KR�9����9�0�(��ԕ+�$�M	s*�O?~�fv=�jU�(����E�$]c�[(:�'�\�F�οS��T�2���<}u
-�R��[C�=u������㩚�A��wO�޿�������R0�]�kdg�?&|kD��K |�3�z����ۨ��~��m� ��(���
˼���F�ˉ�g�����i�}�����S�
ى�"Y�ˣ��ߓ?�Df�����z;�rUG�.0�����jt�?X:�Lڭq��˝����b�*��C�Ρ��NG܄�iP���=�����>��k�֐�ly ?�|����L�+�~;T�lj5f�o��Ö|�X_b����q�����iU�}W��d`����upW��p�몴�Zj��-�~�ڊ�7��-Av�~�zE�b/$K�F�V�����ΐ��^*�'�Tdv+���p��ޘ��N@�=o..d�0 �+{d���}������DG΍���ͭ�uT
&V&o�Ӆ���^�P�&�����P{���Z݋�9����uv^ս_�W�p}a�`��������b̋c���^��ddff&�h�0�0��ں���m�J�\O
b^�\JBf�"*)),��&�I9��T�����v#4M+�� ����,��M���1�ŗUh���+Mi7y��vL�́:U�K
P�+����a����j��D�tiְq�J!d�{҉�Z����uk��BH�ޛ�p����hv�V�����.����!�^s1��#j�wpITelJ����|�L@&?8�2����C~ Vk�Ό;U����;��HzR�=�Pҭ�}�w�:j}]�'��l�0j(H�11C	�j�	Pqkj�J����{�3�'?ٻ�����˴�y���徛�k��%��{�%���_���P��m��M������n�3N�N!���C�.=�����q_�T���O˃i6�p��s?~;]�{�R�������',N�~?ZC�9ȴ��Lx������{9i�Du��K\��.HM~�a0�OF葵�[2���0�f�k_�� ��F�MKq[HX�X�B�fI���ْ�� �0R���Ȏ#��#��O;�ږ'�������_ݝ�ZF��ji7��L�,�?�������t��*��>opӳ�fKl�I�)��f�����^EX��	d��NPu��f�
�5?'@�~���'8
s�,E�ݠ�[k�E���z���S/����z��s��pRB����i׽����߃6Y��!���C/;Z_��%�X6�OQ��OQE�wģ8�"U�I�t���f�:|��g������g$�n�AY(}���@�P��m�ߢg&���Z�-:y2���aۃ�yYC��3lR�޿���V_?��^�r�c6�2�G����H{G_Z���D,q�UXb���'��[�^����hkʨr��(kk[�B�+$�Z��Ϟ2���ݒw�Hc/���]�M��l��p��$�=kGj�Uy:.��i������V5`?��ӀT3+	1+yz7>Cnf���J�uE����؃��֡�v�J����;�<_�}�-���kk���-�\��<	;��Ɓ]Oפ��x���}G��.OI82�D�{�I�#8Ů�k�Y �U�����R5�g���-�w,��0!'
==.#����	_�妺֨�GTU=	��m�8�l�?l0�b�C����g���.�����|*����J0�l�`")�}%i��ݽh�+&e��"!2��&!2��c�}�ID"*�&uz[�;c�K%��ȋ�VSI��5�P>���Eޞz�ڸ���ޱS/x���[�+���x�ض7|���X�I2uEfaĆk������raaa��9��7{�P����<0�{�sB�6�ԕZ�ʣ��
;s���i4����݀O��%`�~�Ђ�D�L�[�X����:��1�e�K��Ho�
��@!�zټ͊�σ�L�)�O|��:�o��;z{?1$��� ���QH�gĳnF��Ֆ����z�1��)������\��v�C3�Q�ìˉT
���T���z���Q�Z]��^����K��^�QB�q����v\1v��|�q0����%+#W���2�ӑ�M�'�!o<��XH�c�; @�?�"�,jbcC�l�q�=/��%o�v��R�Z[S.��:i�I<�\8�st�>�f�+6��'uk�~�"�7�d����WiR`�9
Uq�n'FK`k�uL*�-��[4=�9z�����iik ��p��w��DT�,.|Xoȳ�VVQ1�j0�LmY\;}R���Jp���	��̈t����\�]�B� �o���۔��Xe��/3�Zn�\�������~{
���gq�6]�u9�$�3������7���8� �7*���Iz������Wii%C���xh��녪PRR�:�b���<��",$Ͻ��c��࿷�֒��]�)v�M���L�M�>kv�����[k��K`�<���l.�<��q@�$������%c����yQUn�&�9���?
c����hK��?z9�@#���:���Y��[��2쳰M"��89�4���5���	@��ĘӞ�.�&K���n��.�R����݀V��F�޵B���Z+��WR�T{�n5'���H�n����ӂ�'
*]&��o:�1�4D��ol�ܓ_����\X�
؂<*yK�+sy0D�P���hf|؎΋]υ�O"������E��4
�G�M�`�"o��4~�<m�𻶥��&c<rԞ���	yx1cSΤs�^?�M� N�cҾR�%��&�bh�!��|+�W%o��Ċ�A�B���`"\��;#��g��_`0���Y��:JJWؒ_z3���J�b�9+�}몭\s��44q�<�<����9`�f��d��������h�꓁z_3����q ��A� `��-�x�NZ� ���sH�<���C�=���A��tc��M��ֱ�������Aϖ���Ť�]�jЂ�<cT\lo���勦��(�{���vv�Q��,߾��+ѵ}|y�(,��̌��g��=p����p,t �O����dv�k�r�Så��{���ϔөx��3��$��80�.�]c�
�IU���\�� �wrЦ2o \��ݳ�h�۱<�U��_�.CU{�tN�eTu�}kwwiv�>��=�6�}CB������!�w���O���_gP���$�V�9v��iy��g% �����Y��Q�MNղ�Sh�ƽ=)���;Pj�����#�n��ɴ��e�'�=�'j�����iVV��s�O9H%Sӭ�G�
zN�2E�a͍��n�n/,����BN§`�j�v�:R�P��q�^`�cBޮxH�JJz6�`�����U��k}QA~D^[%(���Ţ�QNCe-)�e��,������)3Z�4A���)�����ހ�Q9V�:W��"�}��zj�>�6G��;X3ť���W����)�ݣ�r�"��C� z����>��L�nIC"��r��du�{�H]��+>�M1v|�sL�W�4�z;]��:?���Y\F�z��ߩ��Q�o�x�{ҵ��"9�����'B>`����H� �/7D��丼��$pGHf����k��CZ'/*���s��[�>{r)>�l�u/���c	�~��h�
���<싽�| ��+�48#y��1����H�S��d������9��Vie)�;d��~C|�Io3����KQ�?{&ո���
XwS:��L�<_O6��f�%5��}���e�\ͮO����������t�������������s��iO�M;�M9AQ��m���V<ݟ�+.	~a�b˳��Թ��ͺ��ע~�T�No�p�bzv�	s��?l�9/���Ae�d���\J�����Ks�����'�i�ro 4$d�+8�Ril�6@�6ޜx{�Kct��JQ2]"vۥI��罗'ʡ�JJz����C@os|u���G2�c��� O�V�8�(��O��,�?��������i�8��&��RP�z�r�|���N�좲�Z�����I��w�[���2���������MrO����n�u�i6}��Q:7��)�Rf�$�(�������f��B����@�?n�A̩�h$�՝u��� ��D�?G{���7c�^0�t9�{Pf�$����(ɱ�ߣ`}G��}A#���NU{}��ma���;W�6����&j�O:��t��">#�^$才�Ç����� �����U���{K���-Bv�^�++�쑄�����G2��d����������x����]�z��y��|����z�^��~�n�z��|�&�n�	3t���1�5X
F��:�ʊU��Z]w㤉��ׁ7:8�A�l��Ħ)s���B|= *���(S�)5L��K�{�j.�ӏ������Y>3�s���؛JcE-����~Qo3wy���@`4�8w�V�n��ߵ�ˠ)�7�����)�-��,��7���УZ�0�P��]fH�Z��ĤOGB�㍍����Juuu@�H������^���?����1�:����������{�P l���C��21���mDZ4�R2�c�T_���r'U:w���|nre��r�*Z�O��:N�Q��.�R\�R*��"�á����l"��?ɾѴkl�{xE?>YN�̌̑,Hs�1��Y�W��uz�6���I̿C�wR�:"��h���v�.�Y�`��Ĥ�l�- S�( �x3�g~�L�#��:�����Z8c�b����'�C�����%�p� �TEm���~�O��X
��@
 �ڥ��4L�-y����g R�t��K`�9`�%ec�E��\�gh���sd�]� ��V��ɯ����.X� ��9�����]=��5D�>����t]���߱��.����|�-�睹����MMW��j'bq�s��Vō=$�H���2���=�.���s=�<H�wmep��������eD2DB��� ��,�h�/��/���|��f8L ��i?����sp(G���+d���E�����
���D�>o��������#�/�p��P�o�0?⣩���e�����ѝ�w��Kγ]3���hXb��뗙�Tʿ��XY�nk��@�NG�+)MA��fhFWhjd��"^��T���ى�i���@'H>��L-�Ő�{$,(�����Y�k��+(��������9Z>}zeii���
:	�A�������!pQ11@�y���vx]U�NI�.�w�ir̇��tO�n�hVd����҈T��֥����ۇ�[��q֓_Cer�2�8ȗ���J:��t***�?�5)���A�%�s���γ�h5�11�6����2�p��g� �ˠ����a��틍-1Ƌ�-��U]���D�n`�y�2��e���q�I�����������e͑)�H�ȆD(��َh�Y¶����Z�^�׋p�Ċr`T��_&LuV<�./���sJ��1E�����D��(��`�s�amړE�,4L�8S�8���r����#��@Ɖ,L��̸?��n� �����IZ�?;H����t��N�#*�N�>��\ %���aEjP��ѷ�m;��R~2J[��V(a��jE�6���L��3ۊN�À��],E�]�T?���?���z�M��t���Uw���j����ը����Ǉ:>���f���=V��5:Jm+�-B׊���/��)o���E��郗%�T��t
\�� $�z�#*��s����bO���u㖇��6��_3�r̦VaajC��"V|����q�	uuw��,r��31=�K�\k��H�s&7���	����EsQ����0���N	:��
�.H�r�X�께p��UņO��y��~��j� ��T�FJ�������X�k�[���Wę�ݼ/��������oO�Ggq��8�L��1��s�����Z��>C������0��[����i�������HA@�R���?�`��Բ��/ǆ���H1 �Y}_}o���(��G	JK���dJ�@�0�����C>��>0,����VP`����'7����n�<G�"x�7u�ʣ�.y`��|p/�����S� &��vw8�OGsdg��
vyXuC�K96m�ޅ{%(}4�;V���9 H���)�#�@Pҡ|���P��������{h셜TF���9���/����{�1�Dl�g>O��v��>'�}޳`�H)�{K�`@��Sr@8_�۷o�B���A譭�wX/񫫠3 ���O���X?���gO/�_��G��.c0U�!�:�=��tm��S�y�<g���3��\��@:�&*hiYH-y�"��뜡����K2�;O�	5���!|24� G�邎�,x��0e�����������]��܈9�OI�Y�_{<=b2[�z�}. 	�'Ř(�y�����@�2&Vf��F?w"��g}��#Ihxy�7Q���U���|����z��]��V���;�#-}������y
�����ҝ����/��(��Y��j�@�ͳC�&�].M��EеB
wSJ�,�ISFF^i*0?T`�ghs����t���pqO�0��!k��o�j�X�8��|�����Wn �l����C���F����'�9L�=>�À�y5��~�%Z���j��rmn��?�9u�T飒����d�>(~55QA23���f�eq�f����c�HY���[�]���o`�cx�[�������x�sV����:�Toan����^���(D��	kc��I�+�i�
:���e��S}��a�߾���Qκ�du�r$bS�w�CUaӽ�^��j ��o�;�&s�ҦL�E��\n]'������k;�&��mqqq��|�f���Κ�׮�KI9��8I�'�Y�?<�h�:����*����W ��mYY�!oj�� ?+�ٷ���)S4ظ���e@@�YR��@:r��1� qdnsI����%G-�����TW�vxz�*N�H���2!/��e�C9*��n�̨���\��o_��dk��L���)���ze+�ƭ���Έm��s������?�����(���L��O�?~�n�	{�
et �Q6���޴��9/���'���B��A��y�noo���B��LrJ;�@��!�����؆�M�����	�{6����D��G
�Ϸ����J�k'�sMinj
��/�Л+)�N\l���!�"����<���!7)fcCX����,@����S��1%7~��↳G(X�_��U���f[���²�.8b�Y���@.i�\[4܀=������2){��>&��Z��EEٮ9��s���p��s��n�a��-�dR��ӿ����gv�˟��E���Y$��r�L���|}�**�D���7&4�u��^��Qʊs�����6���_�;��.i�\�$�ɕ�_��NOO�9a��@���M	ـqS�h���V�89��H�W��=������u�J[�/��G��Xn�?Y��g�X���_�[xV)�}@􆷵�!|������!�:l�6(=�Ur�O=�x�N(+�@}
�6N�am���3Y%=K�s�熬J�f������F(C��Kե�L5`���Y�V�=!w�	�����ɻQ��_��?�Q0y�����4�W�ݸ�z�\k�Kd7�E�wnu���8�{e)�#KJn�]),����;B���:��s�HQN1*丢�b��*Љ�/��&�&m��7�"'�j����!�b��߁�����w�o�鲇ؕ�%K�bOU�ggy �1�=rx^�Z	���f+������.�-�"���m��w��BC[��=E

0k�캟����}�����,8j��-l0�G��5��Y��h�	��)-�P���bL�ܹ��w���bw������"G��1�8=�����)�Db��{��
(�ܘ��g�2��+qW��h���� ^�ҒΛޅ"Y��$��Ç�iԽ�ː���TR�%WWW��Z���Z�FG_� Q�,�!\�9��OZ�x���Z��v4.���f�y5z����{d>Ϲz�%�X�Cك�kq#)q�!gu�m	B:p�l���x���4P��-�ꅚ=%�xע���OꌡD@�#E	�Qv�O��������x��.����l���ɉ��f~��D3���P�j똚�jk�l�*9y�b��<oj��Ѓ���Ҭ�g)S���! �0�}�h&�����F|�O��z~���<��sl[KGx���5F��Up�+�5�7o��¨U��Ռ���@]X�<5/`�8)r<�7�B��|��.��'�:?Y�}�u:�%;�� ���@��O�~�6�K�!��J�i�D*7��t��uZ��˅
?�'�}�ś	TT�l\Vpێ�2L�	�7�4ܜ��n���;���ə�z��I1�4���H<h��4�XQ�xQ&�W�T�����KP�G������ӱ�F�}ij�E/l?�XU���$
�LYF~4+9"�m����ש�C���a'��0���0�e,��R�@�4�`)@ɾ�E�d���'9�|�h0��������øn��:P�����5���%;/�oM=ܽ�\��^�Z���	ʼ��pq�2�{�;?o������d-䟋B����%qiX-&�D�; �͓C��=�$��xr�}^j�5&ff�-�^?�����)��Y��r�T|P�Ql��O�K�(�ݿ��'��Н�V6�μB<�n���W"r���=VA�yC/x��W���a���9/�)+k����oғ��	j�
y�	���Ŷ��^L��(��`���o��6��rx#-Sje;�(���/4�6���\������I�tOL����HJ>il���D��AN��QEy�\\\�R����:���C@ְ3��U�1�8�3���&U#��S"�]��<ćG�Ľͺ�Q[88�B�s�ѱ���j+v�{g	2���m�uHȥ<�o��{{�Z�e��I�$ht~�wA�]��z"m>u���1�$�rݸ�����Ѕ�̡�;ZP<L̄������f㈿������_Q9�x叕��]�h	��Э #����o��gM�>��S�#-}�8���:�{su�P�К��ܸ�Ljo��8*Zu֫��g��1RN�yv�|�ghx�B�^oz�w�{2���i��%s����*=�����\���c��<(a �A�!��=��/���x�0yP���fi�(#S,R~)�	����{��A�c{9���xP�/xe%���A6���>f���%~��I�U�K+��M�J:�!�I�����z�LHXCO�/Z�9�V}%Y����������}y�.�cඉ��oK��G;w9��y�fd����\LA�k%ā|!**��4:kx�̄;EE�A�ϷI�#�Y�� �i	}_�v#VTx����g��HZ`�@���G����J��ϟa�9 �̮a��z�����W������h��M~*�S=/��	5�<y�2Ug�N�,�C��vB�5���w��(��*�U0|�pʯ������w�
>�ss����N-���hW��[{�sp|�����6@�d�tKg��E{��Ւ#^���<�m������{�A;;_QU��4�$ޜ����aw�:&��z�êo��$*�E���_��L�����HP���&�!ߑ!��Z�*��aO\�ґe��k�"��'�G��\~���^���G#yR�x�ī�3�8��S�Hz��R�a��Bj�H�O��E��~�T�K�Ջ���>h I���B����9�w(��x��'������E�؝�
���:)t���	�s���D�+?��f��IJ��cl��V�� �^\ģ��V���ua�����_T=�
��l�Ƌ���0�|.ךxv&�Ńx���r����t���P'����&t�8�������'� ��)q_���KA�'��	�̄���D��P&��1�����Y.01�$� ����X�T��@�OZ���@�ƂB^��	��B�99n�Ԏ�2��hDs��A5����,,����~w���-$�� �蠂�w��K��.x��?����=E��wx8��TTJ�xW@R���5�l[KT��ݦº�����F^��Ew"�oP����^T��L���?;���/��q�ܛ����B^&W�T�IO!�uś�%��4z~R�@��
��l���Y����<VHA�u���_�{��YJ\v��EɦS��TgζbW���:Y����*j�`�����nH�R��Ֆ߸K�ᠽ(ݧ�����Hԩ�m�{t$��m��������I�-�?wvh�%|2���Q'�ez����	��4�d�֯��p	0.P[�c�XR��Pyue,Ql�vC3Eo_JhB�j*�{���s&��G�O�~9��w�`6��UVH��a��<w���G>F����:E���Vx���FY�03��R�֖p�^���b������)7�nF���G�k���#��#�e:;7A�0��n�ʌ�+�������K�Mh������6KJ�&W��Ս��@�R}�̮ޘ�|��8[��m�QW�;��/�7P�j�R��1�-���t���'�7,ͷ��PlZ�Џ)r��~�>ˊ.����/2ά�M	7ZA�+W�\�E����=��0ZͮRSR��R։"F�JbM��.\�"q���4�s=we�z�&�����q�řĦ��y~���aG�*��8h��٩�oG#c��7u��?�(}����f�ۺ''� �$U�v��&����yNr{D�!NN?ad�?�Q��CT��������φ<w[[�n/h��@]t�7W������[^�T&���1C�t(�t��n��w�束�N�p=���d�4��iK�Á�����Ev��]@�鹽nA�gٚ�GLb�6�4[��9��&~��u}��p%^-�����N�q	�X����`e�V#������o���W`��ga�����[��geq���<4��\d��	Vnn���6��wh�`�`�y�� ��*����B��,=��,�r4���r���b����s��>��XҋI�Ƨ��G�� ��x#��9մ��+��h�N,DCHo�wB�n���4�-���������=yش��qh�;d�o$I���c�x��t�dE����j���E�:��TA��^ ��+���-O by�RI:F���a�Z�|�:�;�4����)ǯ�z�����p�q����PQE61�6y5�b0������Ǹ�:낤�ʭ�,\�8����Q'!�8�K�l�
h>��N��F��8��vu�<�quv������.G���Ø]��Գ�'
G�Eu ���DD'�o�>:�y|�ʚ�g_]S�����Vi���VWwwMuuDM͝o��5��fA�T�뤯�()��/н9��C��y2�G�����h�D�p�e�?0+�H��dH� ��q���P��0����G󾚽���wY�x/�s��Wز�ڗ���;�^���m�Y *o_>`��>����0�Ɨ���汍&���i�ts�����<�
����\t��*{>鵴�G�Y"���������z�k�>� ��8ƫ~�q��x�B�U�:��[�K��"{��MZfO��w�݋<<�
��Q��Qо��uLO���c�Ѫ@�;���s�I���+2��ױ``!��(�/4�8�R .֦�x�$�����b���̜��P���Vl����i�j[*������EZ�55
�H���r��^�ٻ��载A�T�Y��Q�zE3�m����!�3��o"���2��2@C�@R�K?��B�� r�_�;�����H;;j�ܭOn�:�_���!�G::��\_�20�ii�Q����b����`z�ID��&��g�	^��\4�ZOC�wG&�$O�5 ����� ��$B��a���m"hl�r�jn��T�����?� p��ws�AyGG6�Jd8U�x�Q�|q����XQ1�1*Yl����s�.p[�����Z�8�`x�ocZ��J�f�f�}���h:65�e(�	}���Tͺ�N��=��e�R����bȚ�~�i����Qi��ʗ��
�����+�́%��d]óm@"����H���rw���Iq	�2Y+��K��
EYRF��{5~�^�+��{�s���j�x���;��"�bG�X\%���%g�Z���h�za;�>������+����F�
]2Ck��OשB�����d�၀шB�8�!0,��B}�]����.������ʇ�C[^��[�_��(���ߖ9�*�-EC��Q++�H��<'�WQ�*%����
t��(�?�:	�*:9�`u"s�\K"�kqQ�1��9���}�]��ZKׂ��d��ß�y�������먃o�_Zg*]P V�v�gz�u�<���w���yh���2a�G��<Y}���lt��Z�x�~��*�>̇A����:�{l�AJ���61��{l�?x{��$�Fz�U@����ʧ$��۬eͫ1���4,Nva׆ �v�5h;=&��tИY[�c�t��@݊���T��ɓ,J^k_\P&��Z��׬���q?�&���%���?�#%��	͝L֣Ňn����\wuo�5�E]U"���ż9��LIDe�>���~�)M2Whk��%@X� ye���;Z!��N(�2�\�����p�{#�%�0WUt�̌Q)�B�dk�X���[�Fme�H�����A:��?��J�q��� $Oͯa3��l��ͽ~N��������Vw�t�1�r~)�����b�N|��cc�Z..�:��4x�0��蹎�<��uV�aa�noϟ��QR�����ܼ�%� }TZZϵ	$:�P� �9	 D�R���0���v����~���knS;��b��]|�������1a�d7��Cc|��R4Ԃ����G��򱧨e�y%0��d���bç�m
�-��������&z7K c�4b���3�H*8ӡ��r����Q7�+W�FTW� S���q�/n�|2����,��������q� �yFF�ی�q�y�z���.�Жu��#�����/��<��V̝��<�>��)�@��0Q%�0%�{��i��w���I��aj�g؇��̢�f���v�:�ƴ��;'�Ko-��.��/e�#'3���TC�
�\���Z>���1*��c��9�?�
�Nf/N|�2��Z�x��tR$v�'��EM�.-�9��Ң\7��CŁ��b�!A"@��KM�������?y2���j��]f!���DD����X4��a�J%W&��G@�1r!N�2;
LU�.z��v��OX��2�j�+��jddb�Ax�[ª�|}W7�TX��Q��Jx���E��x@�a��7�[l�M@�k���1	-x���Qҏ�^A��g� ���[��4u	>9U�?��oX�o�x����Q9��4u^6����	\����9��PK�,s��8��B3�]��Һ�e��Y�0ց�TnS�"�ؔ������q|-���'�/J���6]�&@��[$�sf�	JЌ@F��]��� L������akg�R*4�5���	�#�Y ^ �D��tg��)q�"P�����u�q/��u`�yp�g�����`�+���ˏ`Dި_�L�����P��慙Y�c���%P�#5Q���Dًh������h���Λs~�_GA2R����p]�OrC͞��tdk������ݦ�\Dkjj�����1�VϞ5V�<y�����L��-M�LbjjS���h����cq�� H. !T5���ڄ5@	���|=��M��� eحS/KI���e|?����t��WG>Ua�z$Q��Lͫ����&�Zf� ���F*�S�J�ms�oǈ�k3FB=����U��0 ĺ�~�Wq����>G���d(�����>%x~�>�	�L�&Y�
�� Y�#5��0tJ�/���._B"�����QR�5��}��vu6��i�g�-���'4�"��dXnecCr(Z���#��6?�U�	�b���`����^��i�S�$��NQ�M<�BS{b���t���?.����,�٫"��\�7�p��	rl�5�I��_�H� u���{��T > gi�l\_�܀<V�� �i@�h@�h~��P�Λ�� 6/f�%�%��6�w��VD_#c�
8�NM�,h�s	bN�t�-Q==7� j��;]J�ƢY$�����T���,���u]�a�� d޹��nm;U�=1!�G�����0H�gte��Md�,)9).-=���b�rH:U�ݺ��_��>{EaEA:�f��glf&��X��ơn���^�!a������y4IGŻ��+]�/>a���[=���/ŏ�b!���B�ZOL�Q|%���*��CHJ0_�J�h�w�UQ�2E�XBF��9�ZN:o���h���ޅ�߿��HV�k�OM�y���}42k&�F��ٔ귃2P�DB �Ld��˄�In�J4@�ҦU�^625���P��<(+������6� �b-�<|}���s_7��IZ����,?��c���^P����^��TvX۔�/�o�o��_���>~�B�`rn��N��h�6���� �#�w�U�Q����' h.�U�5*:Xri�� ãY=��N	Y^�(��#R� Y�Ȉq}�*� WXH��,�� l���&
�a "f��`��� ��z��`3���o߾Ex�֕M ��������_��q%�yO<y��Բ�] 2@��j�����a++��s�Y����m@y9ڊ�
tD����sZ�a9uH(H��Ľ��OzEi�y�h�b�c�Z!��u�j��}&�Ӡ�uD��Ec*1�'�E�Y�"fXo��r��R��ffe9;����_
��EsF��0c0���k�W�Z�@F]P SSS
�"p��j�7PPL,�Q��$�@>�yKH$�I�u����7�t7����￢���X�B�$���>{�_ݣ��C"����P��Y�#��J�Tu*B��i� %�1n��=Rj�'�@��5![c���|.���E�V�Qˋv��5_U��Q�\�ʚ[�5���;� �a�r��!�8"�1"��CE�DGWyz{�*p >.�����14k�I��~�%���#�;��������mݸ���&�@���1�VUu�&�]D{o�B������}vv�m�)f�^�\܍�zg4��a�e�|���b��������ݥ�*9��s�Aa��!*��z�
�J����`7o*x���yW�-� �K�hBh(�m�{es �#�{�~�P#��:K(r�3�E�
QE��B�U
�0<J;�������3�=W�{p��]�����Fr���K**H����ﴶ122
���G�A����Xb��5ו�ݮ��5wZj��[[��P�;HIE���� 8OVO*��à�����q.2E��ꌅ|p��>�jS�Y��3dv�\�3y$�%/�p���-P�~Q[)�z��ǘ�& 5��ԯw�n4���7��.��2��\�D�ݯik�{f~g�A���M�AC�$����Y>{��qٽ��f��v��-�v)G��{�������M�G8[[S��g�O�24,SZzG�u>���b��7EԜ^`!�:..�5Ů���-d�R�Qb�u�4b*+t����a���@:(Q��A�1��)b�/{?����¸N뚒�m-6�\������a�	��Ɔ��g|>~bwx]�]J����K�NDq�u�\Hb�x��\jG�� ��X_X~��X�߮c�J��`#*����n��h�WJ����d+Ɋ�N:0
�x�b "%�졻���T�7C~/�)ll4�Ѕ��s�ܙ)rd�z���"0X��|��Q4�~1
@�wAӨxZ.��< ��� ?�Wq����+$s!�@��{��l.���U䢸�$�����d�a�H�I4�l ���U_I}���%a/%�d �������xibn��t��g���=�Z������l��[�Aosr��n/�nA�p���u{�y�����-�э�h���\��5��B����/�y����4�{��&��V�9>�$-�8	p�� X�Y�{C�z�.5!@!OBd�/P0$���:�������'���b�}A�l4���4���v�`H�{��9�7[� ��T�� 1Y��rfX�D��8�9�o� ������1�R�(+;zo�7մ#��'�d����Ҡ�y7����ܺե9DHS�d���b.���&?+�$�sJ�;�g�
����jj�hCZZ*���ڀB��H\  ��\��?�=����z��z��b2 c��k�'�]E�C����dH��� �ygY3�0œ�v���hp �ᢈ���e���g�.��+�CENy����e�LJ۠�*�|��ue������!�)��Z3�і�>أ/���8)�˂7߾�W����8\X-+�,8�
�����X`��/6�T�SҎ�x⌌�#']Q�X�.ba���?���0�ǻ�&��3O����
��)U��SJ��ӝܮ<w��ڢޱԑGB�(Y�h<T�<$̪�]��oc='���䩔��~��6�",����H�{)O?��=�'��+�ͬ�Vl���u&@̓�-.^H��xp�?��B0�Z2[���ʛؕ������c�8R7�A�]�I2�J.��
'�G�T�YԎ%���'�hs�q���32"�
���;�5?Y��"��Ġ�T�d����{|; ���]�L=(��7�/���7�L�t��i�NO��7(;z�Cf�y��s Aк���L�t"f6TA�����2�E*����i7T<ծBa7�:���hq��龶��ћW��؆�nˌ8�wD��߄O�;ՇyeT(	Kx������k����_�8��Do��M��������Wb��?����;�vS�R6M�(,�C.�kp'��?�.�ך5���[+���֣#aqf�9�z�M*\!'77�,���S�-&�K�C����d���OH�6���>��b^����zǦFq����C��_��R�s��f�A2��+T�d����| ��dfib�����l��D@�dr�,���]�Z��W�9Z5����Gr?m�t���P�A��{e�Nkr���Zh����o�H<*���_�Aߘ�l�*���A  X����|�'��u����}D;�Ho��j��]��<�r[<�@MKK�M�/W�>/� �3���_��6]����g��D4(�����A�(�J=i�a���^�?e���,�a���~MS8σd��������Ө7��'("PS�ޡ'�q_A��p�,w�����<���]V 	!i����A����5��X�4ܠ��o��%�РC��ڪK�>o��	jb�;����M�ȺQ&W�&�����m�K�擗�����bT$��q++�?���^~A_�D�����}A��2�Vv��U6L�!�9g�Z�|9YX��yR��z��ˇ�::b�d�_.���iॿ��p�<�H���{�w��S@�:���.+�v;M,�~�\Nظ�0�s$��!��UN���&��u}�E�=�8HRM�U��B4�!w �uFrR2����o�G e_X��=!��6�V��Z��{�H)+��rzZ�իi��?�Ԉ����q%\�%�]$edځL� �[B�A����p�d��������r�{�Nf���e�.I��hL����G�I(��j���>���1�MBA�_̄����F�T]���bE1Ȥ�q��>gı�ˈ�7\+ڨO���@��[R�_�z�r<�w�sUmN���Ag��|^�:- ���d��B7�>O�?UI��X9��;�Ź�t������
:1y�[Vf�=�/��q�n�r,ad�+�����Z�������$�m���D{���Y�˷�_C[�|6.|� �d��޼�K�	�&n[cK����3.(�
h?`9�t.P��*Ε<�,��x�`ÿ|��,�^y��P5�GN���s�Ms�����A�7ڡ�OZի�p/e���)�a2c>��3V���j\�:q!H�:E�埰V8-�� � ��z���'��d��E]uu�}��Z�~��h:t�Y��Xbjj�Q��e�33w٩}�y��b[�˿��<}z�P�,+ͩ�]%�C�k�76����zl�V��:��� �����ꇦ��Ŧ߶�=8����j�A��Ukv��
ex�)�<���]��n,U���
i�@V�Fӆ�sv%c�{���,E�|H�x6��)�l����( ��!�#�ҟ���D��n��>�<a�v���7�Q����w���2�;h#=�[�?�-��h�*�K�������T�7���\�Z}}}�L���6����1�6�KGǫy�%G^�/ww�A�C��[�gϨ�,K���쏏�x��!Si�[�q���E��oH3����X
Fh��j�A�k��є��~{Mc,�<�<AE�|ԟT���/7�l�'��i�d6���n�]�Do5M��L���?�ȉQ�y���wx�|d�}�Hd�\�]�� �ey����*��y^Z��4��b��]�%�e��Q)����aL���{�SY?�5�B2+9���w���}�إ2u��Ʊ��V�=�����z��Ւ_��6m��.m�sq������l@楥� U�Y*�WW�/. ��W)�5p�鱥�mBV�۝���d�F����.3T�׽�IE�(������7��|��D"GE�.����xɫ�Wc�ZO�Y��%@;H��̀����R;Q������Ap�
�&&7@u>8��`e�G���쨏4��pZx��Z��e������P R-�ˏa=��RL��kC�`�Gp��b��R|������̏3��-+�(f��VV�=��11�V;�
mڥ�NA7�B���8(1`�@�-7���jRl~�F�&_�R����R`'�O��vE��	�AL�E5����� � �F\��(M��q��7A���f�`��DL?a���]���r���Ce��ޅ����؞��饋��,��g�8�_ �_�я:-�����[�>�4�ǀ�%<{aw����e���Mc�2 � �t�����_�ܹ���zw?�;�;���T�k�QiDx��+޿ק����ո�|��L쐀W���-��b�����gg2�_��
��u!U�z�7���hv�~��q�O����+�~V=Qs*+.�:R�R��t�������CP�+�/埇�;��g]c�+�l3�-��6�w,�Ot�.�$P�77J�Mp��YT`Ra���!SԾn�졁��0�t�\��g��\�Lߵ�*���g�hb�l���x��j�!������ޞoU0?7�2NS]y-َ�oc:����d��������gR,��9�-lm����_�n��w�1p���	1��Y47Z��sjj��P3�֨���VKojf���_��1��[ʠ�a#���,�J�!�Z�X�꣊!���"��Gʈ��S��e�7����*���KM�����b�kh�����i�/3%eJ���>��ۀ���{Ǖ�шh7��� ��M��8�L�Ԕu��<'j���}���L�G��D���ٶ����/��?��O>��W^]_�=U�R�]պ �v&.����W��������bm��=� H	�i)�s�0"���~�=��^�2vqu�HU�ՁFuZ���{�i>��_^�p�a������-�5�T%*��5_$�|��[��px��[gj��k�`���!*3޼�H����2��тJPE �3޾�9J�r��˂��0/(�<%�ϛC�
p~���^6���:�\�L�eM9l�n��H����>A{+7����QT��F��l\�����h�h kfN�*���^��?''E����y"
����Lk�V��~	9-�4:�3�B$�h� ��Iz3C�;q`���
@��}�l���C��b`)�'Εչ^=���2y�.��v@�7�B���*%���D"�k����EN��n���^h <y�U�X�Q�ܢ�Dux�44T�N�6�,�Kf�eB�pA ���yՆ?9���p�0F�"�pf�;�
:w��\����UX�,Z��2��x�d���|] ���?;y��{?@hC�)⿺$�%���C��ޮ��O
Q9ߓ��͔���Q~��dw�-!)a���:h )촮�X�	=>�� B�Y_��]78c�O����Ԥ�Lv�"~��͸ny�#�\�ɔ_�is��oQ��^R�%�+���/����GT��/� �ɇ��P%g}!7��A�`�V�K��N�P*^��O�i)/CL�-$�FM�ݹ5<8�Ü���n@U,AJVS[{��-��J���
�D�9�}�v�vǁ0�Q�H��5)��\_'� p�\J0��=Ϭ)q(��
�{�@�$@ہ�8)���d�	�����9P8%e�F�59��w�G!�����������v�|ȇ9C���� w�FS!R��1
������tt�*�����옟o~��Xˇ�Hˊ�n3)���)v���d���vw4	wv�Ǭe�K���z�162̿���ՙw�q�P(h���̮.�������@v��k��cuc)�^���<9�~L�o �(�P�'����؋R��X0[��5A���\�����2Kо�L٨����6O�5W�%r��Q��w�A�e<�rswV��ꋲ|����b` ���y�t��i��G2��R2����\��E��<�:���1�>�L�j�x>�x���s��sCFN� �}�q��G@6�5�����	{�u熄�S�v����VW�X�m�{2 �`mk�T2k�f�F�+��"B}ȁx{��UÃ�Cd��� dq�Z��/q��:�q�A�S���t�޸B Τ��s"�29�:!-d�
,}�u�7Ksuo��̙f�����0��S#/������'��H���
���xi��	d�z��X[�0t���<���12�����1D����M(��6p �Qm
������&S��e��a�yXN`����s��&AJ����L���Vf��W#�cВ���|i)hkt������Nn˟�o�G~N/d���9=O���Z��^�\ĘY�W��t�r ^��W�A��/:9�:���\P�}�D���m@�Y$o ␉��7s�c��� d	j�&U�O������,�Y�C>�]� �?��RSS��=qIX�犘��5᳏��g�C����ie,0/S��-�w�0�F�EC���О�o��o�UO�&�;)t�6���.�΢,.�sm�73�O�ې��'#��M��1��sUv�gb���@��;�����zpy7���ȫ��6h�1;!zPR鴂�΄dBH�����&���	-��K�V��_J[�Q�d�E�o���(��-�5A-�->�5!kO{�Z���/4���/t��d�ok�,h?��������Vܿ�p��J�^�zk�E��[[��������>D.
�fFF��!/��*Y��ch�Z���GI@���|3a��ܜS�il����>��g������&���hY��>)������34N;�U)�:�V��v[>�ܾ�HK߀�iS�7�-{X�iH����\�@�8K��ѡ��7)��Ҁ	�}7AN]���b������V�F�K���Ž{�z:-�����X[_�1���kfF�PwEK��/��U�8[��OQP >ǚEq��H�ԅ�9��I���X
}���D��d>" �1J�m�0��@���;������uR2�6���Ҕ}[�йq�g��29td�@�����9D��nSn���1�<�Y;%�(�n�	�b��;�q����̜N�g�eN���!`X�R����ѳ2����ii/��V��5�C��y�՛_)���H|�v�ʠ(��f�*�ץ]�E��w�h�0	�<$2U,h[��Y�=���,+�=zKԕ|�V|�妩��=��ɵ=��n��+*�*4�9�̄��o�Ǎ�ߑ�&���i�+��v�}�]��Ɔ睕���nϥ~�OO�����3̄�Q�\}w<����$Tv������QfF���{d&3�C:!������qp̬����~�����qz���z]�s��uߗA*Î_S�2�͝V)��s :G���	Co; ��x���ڸ�� �ǫ�w��y�H'�N�-E�с�#�-�*K�z�=�sʞ���s��N����"X��MOs��U��%YA�
����-��?�9�@׏b섳�:��!��Y�h��{��.V)U���>��T��˭����B�J�	�^���E�_�V�e|�W��=�����G; ��'-䵯�r����.!�3k�r��������Y�vt̼��R��y������/��,vq�{�sT�_CDY�a���è���HVF�����DD� e&`(Pd4$���n``�^W�����Xoq)�*���,+G��wO�D 
Ϝ�FZ+20 ��|h�CS{�G��%��?��|��P�H`��v07�����e�`��y�q�z���<* x|-j'����<��aWWW`�0�78s\*G]%�\�3]%ze~�T�ԉ�f��5��WG�W�z4�.�w7cZA�����c<�Mp��b���9��U(��N�b���������,���/2����?���"�l,�O �L��C ��(��T5&�z��$01����$��Lֹ�(��z:���>�����O��+&;^���'t�d�hbPӗ�6G
�d����H�E���N~�%�<���K����ڳF�s������݅_�A� �E�3�c٢�ed�����[ncS .�ۡH�`�F��D�yD��,X���@�����Ig��=�@�d��߆,�ѯ
4l��6�0v�G��:�ׯ%�uӳ�Z��ǿ�ml�����=��4+���4Ӡ_�r.�{ֹ.�r,��Q�Mi���D���8�VO`�������d)��JM�;��ݯ�W����h|��<3��o�Wֽ���a� �1E�ܼN9\N��0=6�(�����WE/4��]/�]	���f��Oc����p*�.Kʚ�Z��;J)f�>5�jl5|��s��p�mb�sJ@�s��yO(��/�qwR~"O��ʵ��t���I0[�����N�M��B�EDkɩp����j��;lji�
j��z��eceDZ�ԭ�Z6�$�t�{�\�Mu�Wl�^�{x���p#�cq��JI'�������A�2�<Ԣ�$��nݐ>ZIʘ���]n���k�*���ª+��S��CC�f���M���߽k������������#�1`��w�F|-9d)��k�kR��~ڻ�]Ž,w����F�S��C��q������Q�S5��� �k�'�e��hnȾ�a�"��E���'�o�k�����=�sR�a�Z�ǥ���b�g  ���mY��͡� ]��s����p=�O��+��C##�h�FJ4�N�s�K��'���:�4�u�me�DV�7�Ȕ�0�C����@	�������֒�Q5O!ͭ�?,K�n�9e:(�jE)��D�nLq�g�J���q�m��|�|�/����S���/�#a��;W1<:j9;�hE5}>s�>u��oJ��Hx�M�%	��Y
�]_�VY��ATy��8d�]���ZT���sV*���c����\��(�y��y�!x5�;��<�_�+&0HeW��y\vF[
�'^�&Y���ϫgߌ�O�'�Ϗ�U������Ĵ��F
]�W3�Ǥut�b��)_�'@�U��:�4퀽����Z�D�$9t�HʣK@����5�rNE����-7��.jj�VnF?W��2^�����Y��2�v���c�r��e���~:�\�6.��NA���|��٘;��c\�Z�z��AHh��7r���tj�Y�s�.��:�/��#�n���Z�� ���V����=&2_)P��뷉�!��C¤ �b������}'�Jy~�����*?�VTN:n�>���C��8~�%C�)����(oK,�������G
;�F�����%%J�����D���R z���R������-5E@�;H�+FHD���GG�a*-}6����a�`����P3Ƕ����UT�Dw��_�φ�$��x�p��,��x�Ĕ���vg��;/>��`۠��>��Q��\ZUh���w=;�غP��Cj)����w�����i�_��/��!��b�̒\u*�w,ohh��G��am�<3Z��̌u�<>���W(�jf���%*�!z���������+�^�O�&e����O����h���}R�k��QB���+ޒ+ޝ�������GHG�e��c�m/Q�� �^��ݽ(��%�g�ߙ��K��F��t��i����J�Zb��ƀ�^����j 9s�DJ'S���[�Ul�����;Z�ij@��rБ��7�
��������yyfQ�� d.)����s�����ܰ��u('�����9�r� ��D�=M��wW�ր�C���N���@P����`�������e	��C@&-���F���"���^TD�e�)�_g�'�F�9�ח�|����؃W��i�P������#���]^''d�̢�Z�^����]ԟ�an�OPR�� Ds�������ŏ�O
�O}�1P��j��E�;8\[���^{��iG$\C��/5a<�-˻�J��\ިQE1�{�1�����FC�� �fB��?�Rm��~��U��_�wׂ4<�,-8�Qt2KP[�ݻ���Ǜ�y-��j֮�7D��B�Ot��į��D#jk�Uy���E$'�=T����\�zqZ\����j/+Z?A��<k�n�p�9kr��8��ߝ@�Jw���R�ՌM{JL{�M��O���v����J'����is�\��������ݪ�rrbl)T�����;��=�<�ۨ�q�).k| ~����(!��E��=�����Ef�뛘���/7h��}A"��եb���j��'X�(D�:~-2��o��[v����"q�ؙ)�r��I.#��{}}���O��3^���B�~ �KV�&���V�y�0�upw�F � ��+�N�����]^����7#�`JE5�� ��W�KV��\l"^�Aj���r�ו2���b���z�� `�̤M/r���pE�4�j�U/����>a]���6[f:;��ͤ����KM��o���hxX��������2����9Y�;:����T���=;t{��S�����:��9�ǥ������G��\�] ���I~֭hJ�H)s؃ؙn�ݨD�}P�{�)c��ta������l�ݳ���;��{�AK��Nv�41͘��ഇ�<�>�C̈́�%��Tڝ��]<Ƿ9�6���SL�Mm��e<�z������f%�h���A�^�^pչ�~��$�����aj%�V� h�8�v^����խ����Р����|�.�8��d='~ [)�a
d&�7ʇ�f67M:%� ��XT�}q<m�?�	r���j�w��Ϗp����Oaj*��e��D�}�e����?����|q�~�	oڕҥ�5�_��; ҳ������,#��A{Hsf'����\#� p�L�߇�S�}^��]���{�S�9�,L����#�HX<)?$;�QJl�K���fJ�(�|��x@�,�.��_���뿥&����o�8I[�$�2�5�,��E"���48���t�����!�k�������N�X5�^=�K�b֑���V�G��_��g��yeO��Hr�:ryO�m��6���Y��j��;��|����g���+W���Fi��v�&�����E풒N�!���\k��gb��&�7�ꂃ/dkڎr�OO7.��$��╦rrp�5G %��O�*Zo�d���=�A�s�@�F{Z�}�T���㈏RR��Ώ��jν;_�R	#��t�����%�/����)�d~��fNN��n����>16��M�<; %f..DYd���=�E�����&�#��K��H+'���{C� Z|4�AA5.�S��O��+y�P���Ž{�)\�f�A�d����U���	4n��BJ��Lx���EeX�7�~PAԊ!�5�}���	(+P!�J���R��f/�fD<)$q���]5,����6'k�����л������G7ڞ���x�]	��XB/��3xI�?��V�O}�=��I�W-¶��ϟ-K�q�aI�e؟W,uu�c��g��ޑè�:�oN�Ţ��d?W�po��''u����ޙ��B���!�s���%h��4NL��%Le�w��� �X
|DP�R�6���+�K����g�o��V���$������s���8��m0)+9C���
3|�:@OX��Q�J�	�y9���ޅ�I�l_J�NB�kb�FAƦ���v�܀��~q���,Fߧg6	��b#F�u�B��BW���wg*{�#��H�(��x�9�!q�dnD��|h�݀��e�mtTDuÉ姽��.�������$���tJ���`����uꚩ�Օ�EZ� �O/��4Nt~3y:��K�e�0�	��̐3,���Y]'������S��L��D���Ү���'�
���YY���i��N�ȿ|�Ni�_�",)�8O�]\Kt[���G �:~��{�<�B�9�(�*W����@��Z�)}����Y�|�gKo H%'��Po�Vґ�J�$j�{Jdm�(è�L�˦�T�><a�9닅U��Q�EF����޽[�����m_Mc���S;�qеpܿ{��w�� F7��Q^�Zw�j�I�ϟ��&s��P�k}O{����`�rT�=y��J��'��`�X"PDiC��FEE�}^��[(ޜ�M�	�$�ɺ\��>��A�Fh3�\�����u�ե��.*����3�/UL�[F���T/�� �U씁Wj�bWW�So�.|�7�Y��x�E\Q���1DǞ�U����ɑ���D�Y�$yt�q��r�)t.Te�Rﳿ>�6)�	�y��2��\����V�.zջ�!¹��_C����G��N�u�zc<�ؚ�:B*#~1�D���u�4��ܛ޸���,y&t�v����H ��Ԋ��Fj��UK��M8/��m��z��P�r�f⇶ ���ڳ	���>V����^�z���Pm�U3[��0�����f�7�û�1�(�jNr��G\�fC�͎ �z	C�?�����dZ~������=3#o�am���vu���� A��ϟ��ǜ���l�9�3���751Qc���h�}Ë������.	f��^�WK�X*�r�Slp2Ĳ��4�җv�k��4.|�U�w0���R�	m�s��E����2M�7�<�^��e�xZ��YW��O���������	�	�Z��:7/��M��R@:���ȫ���0/��s�*� ����\�(W�= ��k3��t-�wW�FD�% v6����M#�\;~)�/MHٜ˂[7�Br ��I�G��bݩ���Γ���X44s�wה�|w�q0]��]h����\Z����:`�7�g��Q�y�<a��:�WVW7;`����5�Y]ݸw��1�?�<�\c�T�i��K[������P�RE嵐�}|�V���F�J�`*đ����XRSSe����B��q�=Gy���߻׌J���"$�^�%c��gT�k�Ɯޢ��S�YY9�db�eS��JTy]W/��
�����ꪗ3ˇ��~GQM>�+�g&������!��	�1�/Qy�B���h��'47�xRl)�NMo��5��U#�m,�� O[׏��_��M*�P�S� ���b�f��'������hs�3�Z"_�[H�H�M{z��JD��e��D����K�0����fA1!Q��4?/J�(X"y��"W�כ����8����w��t��s�WK�Ͷ��p���^ꋫv!t�� J����H̀|���g�3��&O��ʪ^�}e��8謋�(��J��w��2������ �m�[��k4������$�~�@m�Eb��:;�^~�M_��m��]���畒j1 �E/�a"���5�����c{�tLB��#9S�A�����MDX��JKd�θm;H��Ꚍ� ��o���BL��\��ۯ���ѵ
=��х��!'�UJ�n�M��%f��#pK�b	3�źF���$�4��EF����j����L7#��_�+��Y��Y��2C�^�23�zU 	��HB�t*jx|\N��������ȋh�Hmz��lQ���d� 01[e�SS[�u�O�ҩh�S��[X��ݞ�6�7Vw�9XA@�5y��������1@&�����,��S�+���1d��S_��W�#1�\�0�� _��#E:Br���Ն���W�Q[�h�P�\sy�C}������d$��2Ԥ�z%z����5%7���
 ^tRUR�����Գ���J�g�J��G��1��
���ۻ[�O�;N��������MM���KM}������V;~�Ș#�nm�2����	��qBE4��c��=��3��bFڅ����,�g��v�2Y[[�"+��W�.w��_r�S��J	3��Y�H�?0V[9QkD�>�l�ܤ�_�����kp8CF-.��YW�����ux����"�T�Wr e�W*�}z4���3�=-�z���0���-�gj�&�aT*:���*^`�;�g��E~�E�1�J�:�$���s������"��A���p��KW�r�ХP�?�,_n0ps��'�F�-�1u�G{N�-U�d��}Y��2����"�춸.4�����,d�+
/��/2�H���-z#�����������4s����4��d�/.u< ՚�9�-ѫd�>��j%�Wv��Jr?]�8D��2��+
׺g7͂N����d�m`j���܄
������@�����á�1�d�`ɉ����Kk|����ϝ�ɀ� @9����9
����f����j��2���_�T��ԍoFΨ�^�<41��%[�M����e��8E�t~�p�H�Đ'1�2c����(���	^����ش
�(��Y'm����@�,�W����$�/6���:��KY�e{!��#f6N�sX���ު��us�4������/l��T���@w�1R�;Ȏ��CI����k�8*+zc�I���Ӵ�U�/��(�a�L�K��b�nii�x�L���q�I��f����_�:�j���W�}M��,�K�u���� 7<�~Kk����Y޽{WS�4K=��S�bvM�?���eS"��π[�	�Nr;��#z]�}y�k�u{����k�Y�,���VF|Q�&5wف*P*���0�Y�#�QGu(�(p,p��ͥ:�$��Q�u�C������sl)@w�T��S���U�1A\W:K+svυ����iW3TŽ? \�q�����g��L��ל;��j��E@�[f�Е�]s��
�@ƕW�W��E��{{{�Tz��ַ�����Ls( #Y>�P�\��Y.f��;xH\ZZI!_92�,�����j����Ο1%So���8̒� ]�I9h:K% �djo  y�*���qH�����̄�?�W��L�������S�M���E��x�����a�[<Xu������,����/�lF�䙡���F�pz��*޷�ٷdԸ�HL���k���� ����#}�)R����|���tu�wP��ѕ���⧾g�8�v
z�Ƞ�%H�ߤ4��Z880���{ׇ��[nVY�o ���J��8^�2�444�^�VX��޺k@ I��6U�� �_{���0)�n��
3x�R�,N�)�}F�Hr�TI���Dھ�W(]�b�XϚ�p��S�Ì|v�נ�Y��� #0�zH�T�H�P�eXɁ^P� 4
{�OPr��T��a�zc@�Vx��P�k���Y#��seďZp��w��#1ji{�S�=�AޓrAz���]�ior������`*�$��w��|Ũ�s*ڸ�~ꏗ��f`U�P���j2����g��kD��@*�8�Rș����H�Iw:YY]y�W�d隴EeAL����AH���.�{4���Y�o��RӞ���>Ɇ��5�{��$�X+e�ue�<Jo��w�w�UDop	����_��n�L��VN�p0�0x�`"/
o�7,ႩD��6�Z��$Mm�&*���:�����7�� G��n��t����l��pBҊ!�������0N�bڪ�1J�BI�o�l�R��{�gǾ��I?>��_��l�w��]]���f]]`G�N�n�}#�Z�8E�23�<�Ia9<�Eˇ�i��U���U"��ݎ�\Z�l� ���QB���z�������X ��
��`ޓ����S<Q11v�����99L!-�R���cb����z�^1���E�s��������=�U�l�\��ϟ�����(���t���r�y��3��~(�phg͜��A�O:�Q
9��]T%��
O���mr�Q�E}��E�m��":�4��B0U�:#@��_�Y�yOB�/��i�^
��� ���u��
�#n{�������/�P$�%QWW���,x������YρϚ��ο�#:[#�W~zpB�2{�C������go/|�6&��m�w/�X�Ei����b{4_�S׹�qlL����-5����cY \0�O_ }��zqQ�TT�w*.v ���.7�vhN������89�K%B��qr%��m?�����0C��8Ӹ�X���F��g=���������) �[���	�$2�j�&(���%!
�b��}	ޏ���~? S���0����B���'c��Ն���\�9��l�Ed�M��B��4��Q��V��9��B��.�Doy~�
8=�M��\ڳ��a��$D��x�W}�������45>'�#�kU���j�I��V J�"oQ7���𦚓ఔ���Q	&��dM�w��Ltʟ��4M�̌<����Lq$^6t�ތ66��3�c���j�
��u���¢w�&�բ��]�v��,@������Xh��-�]��O�c�K�(��&OB�ë ���@�E�j��R��כ�ƺyO��h"sx҆����^�\={Y�T-��5�T�$	�_��wY;�t��o>L�-�9�+O����.gȁ��v�=/*'�<��겊?:�z�uP�&��v�6�4mv�vb�t Pϖ���i�����ʥu͂��1��|�_��I�6ϊu�kjP�L1�����m--3}��	hJ��3�%�s �w�û��kLSAp=	aׂ(�&~��S@��=�����j&�2�.�4��P`00((E�U�Ȳ@KFv l~,�]��,u�n�IP���/̵�f�z6�� �:K+A��)���,���S�C}):g���;�{ar�ߌ�����wU�q���⠒ccjܡ�sB��
�cw2����a����m�d�g����wt�b���1O������y�=~�X���.�E�z:��0A�iW�t���X�UGA��Oxq�u����s�����5��#�@$991���.��R��&Vђ� ɡh�w�#�J	������X����(c����@#j�q���[�:�k5ת�W[k *�."���i���(�2Lb`��1v9�Q{D��=�J��W7}��h[����4���)Æ��Y�$%{@W	���/ kUV�����\;�8�sz�$H�S�M���)a�� n9ӳ�?c��,���a��4�ǭ�/ƤN}��)Y޺����'�f7X��r�ۣ��mIIg���]?�^����ҿ���dT�IY�M���Ʌ��n�C�ǲ����z�&\���C'�������	�"�Ȥl�ϟ�qq�!���甾/@�R�Q�mQ�eW��b��nTc뼆[��_��y�o�`�{-ӫ�s^/��)�X�A�æ��������r�έ˓�c��o�Js���HZV��]����P�X"��� �\q�U:A�3亂��8�����u`I�c�%�T��þU/ɚ]�F���1��ͻ�2��M�{�o�OFWi�N�M���c���rp0�8�@}g��� Â��UJ��R��^�����G�<J��Jɡ�K�rN��Vt�������]��[��JF;-��B�f�KK��UI'������^�Lgw������#:�-�A���4���p���E��#�=y�qs#�V�jƦw��{�p��Q �]��t󼜸uje���|qz���%i��NM�oh9]^+X�M�91��H�J�d4�n����Fδ�J��
5�j�d��K�?�	Ϸ�I{�w����8ch4��!N�F�f���m%#�&�h���%�.t0�.�_^fL�%G��/G{gBA�	�ĉ��G#PE�V���e�/55����F.іBỻ���$�|./i	�ј�;���˳EٵU`RD͓vR�q����	ҹ��('�"���;�	%P�|�g鉰��V��+���+���.� �+5Ռ3��7�{2������?}�/q&��]s�R�!��o�*è�@��@7���p����]�`.}�!�|m�M����7#D����B�C�4W�+ot��,VT	҃��K�����vκ}.qN��KJx1`7�,k�;�ag]1W�5@:~o���o�˝!�#�ց���@'m�:������%P���]c	�+Pk�T����MMh�j�d��;wLE蓭�+,R�/{��\�{i��{�6�{�%�"V782X@Ƶ?����Y��p�H�pNp�5�*���Һ�;�P�*V�9�=���'��z�+���\�{P���FQ��4�W���J��f�8�\���*[�jÍ���RiC�Ld�Y��1��ɔ�'A�h[�q��hԜ\v�؉�J���d|���vSQ����0x����l/I�J�'�� �7���BC˚1�X�=�Ajym-���F|��E�	(k�A�����F��zpdr���R�L�?������S0�q��(��͂t�R� 	�w��v��6*�ͬߦ��c'��RȎ:��˱;mh��
�*�DF��C�̓�^����"[5�+Lp۵t�=�����beu{�j����o�r)��@\�D����T��[�,��>	(~�{�2?2�$hR왨/]H�Iy��O�����V@
cؙ��������yD�G�,N��
�A�u��)@H�n�R�M�35���kE9_RI�R^n�b{kuL�'�h^+tu�+C�0貚�565̗���-R<@߃N~D���6v��Y��A}����u�N��hZ�L�3̋�( A�54�|��;���x����r~�QVY�]5���h-[��IǴ+�� ����'Ag�0Nbt$	(+h�f������-��:���?�	1?H���:��I�Fs%�։�޽�9���y�5�B�<�0���o�l�ۜY�c�1�_������C`�;	v_�d��	�b���:L����N<~fd���h^+��K>~~���1������d��}GU������<�
�0T�А�,���ɑO���a9����5�<�-��39F
i�?�Mf��C\J�D��'���/��7h�/���"NuǄ)��M�gĔ����}��	���MӮM��;��d��II"��K�P�4���'#~"�TJ��Cz�`���]�ڎt�q�tU�,b�>/�jÞ|O��&eD� A���J��c�J��9����1Hd�f�D�vG9�9��@B�F����ꢥ�g�m�/e�bT�ΌD4��|(;?/"}�7'�K�*�>'�O�
��ݭ
ޮY���U�5�]]_�G��u��
���:�hRV.�ǡ����O�I'�IF%�� KJV�*����I��=aq�� �JCC����
�>�vzۿ{�b�$.���ϯ��/x�@n�!z9��"'ϼ��:�|���)����բ_���)�a�aT���:gAm+ek��/��>j-��}�͆L�����Z�EP4h�I*�<3�t�2�7�)�K��?|����)���,4,5r�I�lÒ��.��J'�d��k�/d����A>�ABJ&�(��u���oJ4t>��r�S��-�ۺp`�

��l��Et�\�mcly��OO�+��--��?k`xηI/2>A�*s!�?W����,pd�w ��%��ea;����`��@�_	�����R�z��v0�'�2�g��7 �9@�����}��\t�aI����=4�w�L�Z�)tۭU=%lk$�:giR�r�t����Q��^���� ��~M�?N�J@TM�=P����N���)9�`�2�J�/�E��|_��*�HU��*ް�H����ߜu�=��W���}��K�AH�D�ɓ��O��{��"n�Ѕ6N/f�G��ԍ�\�_AۯC̬2@(��S+
������!㳲
 g�~��ʀ�;A����M���w<�֠y� ����$ؽ͙vJh�ʯ����zƑ���mYIO}��E߆��ҟ>⺊f6�=�B=w��O���Ks�7K�PՆ�'����\�j���lEt�Q\����eۚg���L��K���i-t�u89��o^'gKC���'��QhR��L]>�VI��Q#��s��*����Y���p���]ÊlYod���q2�oQ�=e8�ol�i�������]"kxt�fI7��nm��lF������D�ڴ�F���mKSi�}���rZ�,+�{�� 6���]jm]]���Z�{�Ғ�н���������E1���=����������̓���&����>�8nLQV5��4⿊�ȿ����ڻ��	_������'0��fQF�(l�e�=4`j;�|�2 _�L��\u��V��7�`��?ۙ_5,#���GK��i`>����nK�!S}�
���~��3f�Uuu
�-jjjb�g@Kr�L���N���?t�o��F$��A۞��u̹�����&��X�3�QMe�75=���3ڜ�E����=7�Y4��=<���Ws�򂐑��{��)"{����^:�ׁ���.�K"r��1��O�
�\�U���\F�S�eXU���Ǵ�����sRV����X�ձO�ֈ����I7ޔ+I����D�^��5ⷱ:l4,���q�b˯��-������ӛ��v��f=%ж�}˻�%�r�6�.�2_&�-�JZ4������Y(�%v�4� �5�)ʰs����* ���v d��!���H���_�u򵡎����芵��5�k@@��uk�I����@�O�����a����B/@�0��f�q.r?v���y�L��Ռw��L0��?{�����5DTV�r�'Zb`g����&�uW���Y҆��/����Ra�Ѷ��9tx�� Y�p0��hlP�}0,}�&���}:D��+`�̼H� p��l41𡃀  (�O��8�u�(Zߨ(*J*]>���u�؝k;��Z����jP'���u7��殪ި��>���Q�1���QA�9�ތd�Oہ��[�y�i8�%��g�ԯ�*�˟��*�b�~õ�~v���O��#a���%�~7��^Myt�)���	��h��Z��
�h��rt@�&��<iUO�����K���f�\A��us6���e�r�)����0hG�R��EY�}���
��)�[=n�9�Pr��ۮL=�-�QKS�P/U����������}|Y2�z�4��5�\����jG���S.��э� o�:��ù;}�ޝ �:<$�R���3fWɭ���~�tlmQ�m����{M�]{{$	|�w%���7< �~|��"����薋n��1�7����� EL�h��}utn.�@@:��O���G]]s	V���O�� ;��=w�6��XwO�X��@���3U�=�o0?&��A�r��x@�v[�o�p3�f��bgE&U��$(�TE�"@�E�Ղ�Ńm?~�Sc�x �5_-��HlN"�Ư���tLQB�R��)J2�gv��L���y~����nD��Z�����;q���Div�9Jd)I:ksf+p����131���	Sɳ��Ŭ�9����6��R�����)O2��B#~���{�݊G�k��Y�6��!M-�=�,��/*��n�7�Q��J�t6z⵭p���c�=��ҏι8Gռ�i8T?��J	�ȰVφTpM�>��!�
�<[L�!��>)|�t>�
	��fR�پU�ioU��@��ظ�:Z�b�@�ʦ�����B�,L�K@�RC��H_� F�F`߼�腓�oK�2f�yB�Ԏj��/�w�SJɿ ����9<WD�j��"�镕�|�7fa��^(k�V�/��$%z�|K�	 �DEEo���tY
:��%#�Y߳��"%g�k�s@��=��OO_��K��Hr�"p̀���L�]6)s�d7*���D.��n��&����DD�eZ@G��3V�mK��<˖���~�Y_��C<��P�˺2sXF�i`n_�n/�E��5�~���̤���zh�D�b��������#�2ktڭK�9�Op�+4��^�
���r�B���u����o�ju���a�Bi`e����C�����,�U�=pl��]��b����8�<:��.(%��kk���3ZP��d�Ak��
�Ά����X5KY�������S���;9�C���%^�+6�F��P[�̓�X��� ���j:�׻-�$* ���'�(��e��� r�����B���Լi����Tl��Z(�viD�Mz�\���,ʉP����vtX.�'����Ϡ�����4�r��н� ��w��xJ�E�?;_��č-@{�{���=]Yo�!"�Y�yw���}�o,���1��1��� m3Y�ux��}֡F��u��7q&�����1�FcU���y�kk_�ݾM�u�1q�87����«Ԋ�L,��O���x�2�E�O��PA��EYA��6�6!�r��2��|7��K8iѕdN ε~b�/0uW��ڦ/~ʣ�n����a�I��\�����8�L��f�^��Ȳ���tx��6���1����,��6$ض���D͝.fԀ'!W�/0�xS���bY�[<
$8�a�����سT����fM1�E�2l�������
;K0���B\#���B�`��끈|����
G�{��+B�����O.;��X޼�-sTV�u]�eyt��κRh�ӕ�') �P���r�"T����DD�]�}^�*��l3.�k��Aj�fxH���5�2��J�>�d��=�G�!r�g=̗��E^��~�	�Έ0O�0�ZU��]�M����؊¿���k��\��I.��8Ĥ,�W��pa��EOB!�&�������0kP5~Q�iJ���w� �7�C�����G� ?s���Ɵno��;&L��ǎPo�w 6ؠ���(��G�
;�˩DKh����3~5�zxx�zU��N�M�]~�%���~�*W[�m�JRx܎���F�u��)�k�h��@~�u�qp<f��z�[S�8:y��
 �D/����AZ�/ȺD�
�T+��0�T����9+�V���fP�N���!(�+N�޿��wA�+�b��%Y�Zot4������uN
bC�k9Д��v��[N�q������mTuAٔ�s�����tz#<F	����V�<ޡ�!5F�0���ɹ�vA��o�E/�̂�ɳȸGԢ���˳B�� ��~h)��#%�b������F2"Y�
�1�_��_��w����Sʱ�{�����U	C/�>��^Z��F��e�B�{n=��0h��=<9��ZŃ}KU��|Hr_���P�S�Ǳ� <4w���(��i�>�.��V���1H�4Tx�t`��VX@R�je�;H�t�F��J@���ɓ�Jd}�./�P�3�eRȃD�>ϧfݓ;^�g�8I/s�e#U|	���j��}cbbRi�a�<���)jA�#�OO��^k6��al��璒�}K��SU�V�b���g���7VF�Rari[�R�Ƿ7���lI�>�Ft��J�C��/&�G��׾�<d�;���vb��;����E#�9h[@��Xb�A��3�./I���� T#�����.��'M�@ٚ����#�Ts��ۦ���s�`�K���y>�$P���F�Ӛ�7\�:ʜ�@疞6iH�_�W{�)�L�e��^��j���X憢�s�"�V�X<d[���GlTSӞR���w�� .�%���e@�_k�J��\]���M��J�,��ʱo3�,���H)�?�[|�P��&&!����s5y@f�$�#��U��T�S�X�$�3�䣨���?�}  �EL�N��\�����������9�KA�ޭʲ��
�A��|K�<�v&�t�u rY�j�� Do]Y����ir��(|�_u�I}?�ѭ�CF>pN�]avě���	'.���7���/uJr���TY�L�xf	�db����z�2l�����O:���L�4*5P�Pkg��6oEE]�����X�2+B3+�Q?؜L쬷����S�$44��p �O��	^�@#���ϼs8 Z����&�ս�||J�S[{�[m=�$W�]���5�㣩����@���H���1nZ��H��HyP:��E����jH�	��1'a�c2�K������ t�k�P�\U��U��6�:��#����z�^v�3#fSD2P��7�.�P�?��� ��S;�?C�C��KM}̓B�5:��I�/�|h�jWϝq ��S���@I�{qs�߻��j�����cwL���/��܊Z�����ɧ|4@�^m���>�v�!{���m9���w��w�USJH X�|�A Kޓ��56Q=�H�$��ԙ �0�.�<���]��@L�m䵋�� ��U�3��@mZ�UA���{���eM:��w��XK�Nb_-A�F�X[ձ�����aB�G\�#MC�_�іע����t��<b��|*�;!|�|	��!�\����|��؀VI�)"=<�JCN���P>36�������VB0T��ms�fy�ƹ���9{�Za��8S��V�\�W�zh�Oc���ny�	�ɺkqx�	9���
�sv�H[袡���c�	g�2Sd��&e;%zx��ز�^��t?@��S揫8�k��
h{�ڔ� �$t�0��S�1���.��w �@�
�RO�
�c��4BfP Z!+*26�u�P�[� �����S��¡�m�S8�Y����ָ^,�D���ja�sIŦ�u�_�|�hУ|xCgu+�a�Ȥ!(�I�6���� �kcM��q�S��.�_��r�	���+2q�����9�5n��M���|�����.t��4�oW�J���:��N�9֋wQ���=FY9����5�AAqzŗ�E���u�0��,���sYl1x���P�����I֗�v<4���owU@W��B�Y��պ��w��������Rx���.���7�t����7�:~,��p˭~���!~'[�rĺ��6u�� ���%;A���1��~e���뒜j�'[�<�z$���ɩuk~X7�k�$KGggi���{��9=R��4蘟w^���E��<)N�.�ɯ���LΆ'i w3X�Ʃ�����[xx\�:���/�C�PON�S�\R���y=d/���h 5�U����z�(���R�.�����
HHJ9��t�HI����R" "�0CJ)�w�������r�Yf��>�{?�w��
vk8TV�ʩ���t��ftx�����,�[
N�� } #��$|g�Ĭ���r�c)ly��2�أ��6=��pΔL��m�$�GS�ߋU)��i�)��T$r��[�_$c���eΐ�.��i|����[]��1��.R@g���
BɃK�j��������H�>A�;ff7F�N6�y-�7��X������4��3e���<A�l��Ѯ�� �j��f���o�G�0�_�vLW������Q�V@aK�k�T�|�ᶛ)�@.X&���N���ѡݹ� �6�v!�!�I���-�s��ܩ���k���/j����+5�k��n��Zq����;���ds3G�׽9����+���i��2��o�?
����G}گ��se��= M�o�Z��f?n�����r�o�X��;���{�����H;QX��Ύd[��}���d��pm4�3�����1�J���wʔAZ�;����n>߅<g�S��9z���W��](������8���/-����
G0�8�D�.gqH��m��U�ɰJ�P_�5j�w	�||�T����c"@h��'=!�5%ހm���7�\��b~�����X���a�V���2�QD��JǇ&د%�D�t�A��۫��fF�MY�=�j@}�e�NN��*6nF�8��1S�Ő�d�G�#��ˀ�*�T^/��F�d��<�����8 ��q��Z2���+O呕4\�����O�&������ɶ��:��� ������8:2�-�߬����<�r��9!-@J�mRq�\~B��z
S[��Ӻut�{z��V��:��ٯʘ�;٘ݘ��]{�l��d�����}R��7���B�$���R	)k C�2��8��X$��]�!�C_}��?�'6N7�*[����m�e�P���Y��՟]�����k�g�r�(�j�r��_%.��M
·�Z|��$^0ίR���Q��w�ٽc�R�ó s�����&� �͖��v�[jJ���Y��Z�����)-��T@iV�ܣ��~~Y����>r\j���s��̪�c2�e�c��2�p�n/�O�ڗ�U��M�'�Ky�*==]Q�>�	<ds���n׵��*~T	��ME�$�<j�h)-M�����2������EX��C`�S�o�$� �Fv[&<QT���"��K�<ї�	r��`��\$��f�#D��ߥ���HAV?���\�5k�5V�p�:����E���9I����v�
;���3�������p ���j�����VVV>��L(J�juO�)x-��0�^�KaqH�t$+�9n���r�=Eo�Em%F䌅"��ᴷ�UA�&��tq��#]�z�!ul��U�b1 ߿-퀘~�UBSV�)vl��Y^N�c�JI��߄e��˻�{o56������}Ƥ�[l)����rd���q�d��9q���_x��eh0������D[�1�<�]kt�ѿ��/��l����M}о0C�.���F����
ʣn��W�E���9�[#S�R����َC-i��*����&��O���%V��#JK�����ȫ�4��_���_��Ѝؾ�s����:n�~����l�J_�+Ji#��8Q�;k"&���Xx�^w|�� �o��Q��BP�Hr�c�"n~���AWW�&
��	B{8jobq�/w`}0�����dO��T·�����<<�Nl�U���5ߪ�:�;̴�M�����3��]����:��@Zh��Q9�4��d��*-��q�lj��_f��,���Ϭ����4��ci�=Gk"�u��퍾�Lo�������⌎x���3��_�>��Π� )��u������ҏ˲���� ns�ׄ��t1����-��!q��=��BQ��GGJ@d"3����C!de媡��1����~w�?�h&�&E,��G����m����M@��fM s��Ng�s�:%������ڭ�o<��ee��ml �%�� z~�6�p8"V���h@���[瞯���滈�_��r��� �pk,'�S#����\��!��k@��� xc��L��-���6P���RiiҾРl<����B��4�<匋D:�.���wp�0;��l��f��Ⱥ����EtY/��@�М��h���Ғ��������w����o�w�_A:8ˁ
�F�ffpp�����&|��ƍ�:����r�Y@'�k~�_�[�A�VIhE�];
.����us9]�~c o��q�>�)�D�
����y�)�NMz~��\d�͂o��hph*ڣZ� ���	����z�)<�eS�>=���6L\���C�@���B�I��|\j�u>ݾ�Wh��Ӛ�𒎈 Q�$�M/1� ��B2��Ǒ5���Np�|�XX=�V�k��v򆍈�������J8����щ��=qs2w�p����V1�0�]hx�[�(K�Y��ۨ�ZZx�I���P���{�k�Ѧ�R�ԥ�_o����͚��u�%5��]�h${[
3��/��J䲧&�����bh���@���S�3�:ԉT&��FfOD��C~9J�P�~��^|�D��'k�qqZ�ͫ��̓�1'7�e|hp2�&�4���(��v�m�X;���*�pKKٲZ��o�cPű�����\;��Ԋ��>(��݋�����˥�?�5E�/�+-=\-���=r7��8���I�S�d�}n�>�Wv�����1G������:�c������W���>hj�e0!�}6��8ܾWT���w8F`W(&&�4���B^'�����V�����Mfbjj��9゛��@��$��p�c���M
�QǪ�ue�D9Ą|E~ɠ�G��rn/}��g'D�u��X� �L�w����mo���|�y����.�n'J��r����*m���p.7���FȸJp�O���������C�R�um�u-?������~�#�9��{⵩�~���)"[���"B<ى癿?��zn�)Cc�X㷶 }��k��GT�����s�{����ZU���QG�����\T���W���������Yn�y�U;ق<�7[��fB�AOZf �!-���a��_+���m��X�ҫ��9���<1!�C�
¢��@ s+��su��=��'�z�^�C��Y�CW��	���o}�����ӌ���m4T��Ws*.�y�=�p62}X��<�F|�S������hDt�2�!{|m���}����4�b��|}�[n?��)��%������#�h�<��KҀ��ʨ�'O�eɱ��i�G�fEB�z�����:�"��3j�<Wu>[���)��u�G���{���z|�Jx@�}V�_���U@%�ra�k	/1���̠I��G=��8�ԅ6���w(L���`�bY�x��C��#Wl�=֊��]�A(��k�(�L�RM5��u*�_7���Aw�<��	_{��<�}~������c1��,Yv��l��4t�{���"�j��}��nB��@��2)�JE.��n|��Q�l=�4'Ue�pޘ��ࢢ[H��y�ҪkkÝ`$A����m�W�ۻ�'fm2(�͙��P��x��������OS�%��������0.�9�y��2��t�{�q.ք�q���A%[�ڎW� C�$Xp$b��,j*�{랄Ն?ܬx�I6WMF�i��LQ^�śڗ�V�g���߸���*�:�(EȌ��fE�أ�{�3������4���O=�GK�}��X�����q�8௴������^6�Y_�V�	�u �R�2.i@h5
3����7oȇ�=#o@�z7��@����:ܺ~4bk��5�T~�1��)'��|	&^�XWa^�!?u�1�;��|A ����FB&օΘb8���\t�׀E��N��nP��`�rr�$��*��� �8t�z���|���_��ڛ��_�d�=8c�A��~T(��?��wI)
��d���啕�'�k"�����k�qs��ww_IӚ��·oV?�J��_113����Ԓ>5]i1����v
���q��wu��]��w$B�p)��2`K��	�R	7�=p�cy$~�zl5��)��#^��S����j� �L�M�fb�$L��.�	4�|�;���.�XƜ%�p����Aو�L����Z���a�|��B,)�E��]�����q70������\1s�C�Û�z|ፍWpJn�;�X��������.r[=���S��W���kۼ�8g�w�`�jRX�=��/���#*w>�*p�p�`f_6��v�������.]?^B����բzI2�u��ݽK�DME5,��� / م�]�����r�;�e��L\�u�O(��@>��ө0 TV���1E~u�������dlL�Y�GX��-�\6%]`�q��$s`��L�C�B�B���k����a�����)����]�*�7��v���%� ��ϥ3[x��7e4�7���0�l�o�O�Ă9썑N0h�g�+��--x�ӧbhAҵ5����^��������g����,��ݯT
$'����%500��ev����.+�Z��s�A��N��������C�]?:�d4�p�ꜯ��QDv���Ӏ�T��}�C���#�6�(�^b�����o���vf������/��w�s�zIY(�>sG�;�e�q��q��0��׸,i�,��Xd?��'�v�*^�[I~�1l��a�[�j\ɋ����n|���Q����3�H�K�3U�[HL��5����� T�7l����F�]ֿ�{_G���#�*WR�t�` 6�`��H*"�.�<e�B�Y_�
�}
_�����Q�W���k�-E��W0L�w�@�ݱ��@�pP�k����eQ.7(�o��I�f� 1�ߙ�hVE���B�K{�zx����*yј&C�D�m9\����]�iG`��/�N�e^����S��o�oK���m� �+��4��/=��vln��O��^�z��ys��՟?[��d��=<�V�����!�!.<���|j�@>�zC����4���� ެ�N*��	IP���vc��8���cm�,|�\�R�/%2;�%�D��
E��xa�C�gYM�}Ax|�<����y�5��6�%�>3Hew‸�@���&��)	���A�;Hw�1{X��0�36q%�.�_MB�Ç��@'+~��8- �&@�>�v�UFD��I��6J�%��U5 �J�6�/_�
k &H�-����>����d�O���c�����1���. �CHx_�#��>F��11���ޤT���!145�&ڷ"�����Ąb��bw\�n�����ov0��׷���K�o�[(^��9b`jJ�8<Ħ�7��|:�w�����A��T744L:"��m��&@l6|��ر>�q�Y�H돫���f�JN���F�=��,��G4����x�m��eX�{�qY@|3��o{!_;�g��ϟ[�H��a��� K�ګ%�����rFĲE���}��\,%--_m��2'b�;�~y��'"�'�Nk��^m���22�[����\���(�3o�?�!�ӧO?�I� ��GL4��E@���j��[c�*א��L�|.k� �h��ꬻ����.��O�?�B��,�!�@�NOZ������� �Љ��dk�r8(J����Z���)�rx~{nu�W���B3ZY�!���e?������m ����(;��_��ۼ$����[��������;��8ɫ��"22o�'����G�e��'''�"'0{�<!��_�|IZ����y	S�u��f�����}���.��K]J�)���Jה��J����U1G�٣`�C|"�P�v�<!��o6��{�=�֨�O7fr��5.Q����]ܼ�LN�f��M���r7}e�����Z2&!�^oMY,��A�������6R�[i��B9զ���o��v�i.�ŞtܾlG�*B�2�f���l�?��W#�%�Qj�oi;i�`WU���Y�W�~dk����o̞K�Oe�}5�G-8�����o���̪��U#��W�"���-���"���f��ζ��}(��'(��L2x��8����@��CE�]ŷ�6~;(Ւ*Y���6A�����
���X��e'Zγ_V7L�_B��fW��o*�	�I��u%ف��ٶ��bBB�����1�~)$R$o�fV����%�Y�k���3Su�=��%��T\�rL�����M��.r�R/�'�./_b�@���ӏ�ŵ5���h":::�\9@����%���e�3�-|OĚL+�?�tR����bFōD2�k��J�Ԥ &���_iz�D� �"�<����{{��������b��{���F�&��0����VX�A�XV���8|�4�>�� �rҮON>;G~v�v��P�$Ƴ��8��d�(G_?q����~�J�Z%�n����:̡�4�/*WFӹ�����4��-K�}�?�R�w��V�`{���Tb�׶3ƌ��|",fvw�!�e��
�뻍�4���v�z�j1 �[dr2��$�7OY�q���������ڂ�&^626�y&��1�^����H��1�j��>cv^^p ,*|ိ[���Zi+i����'�[(���m��P���}u���⥦=�qq!y<GT����U9av� �DE����=����^+��2S����&6��^���k��?�����C=�Zޡ%Ξ��Ŧ�h:K�p�Q ���O�ޘoQ��41�O���N����1��
@B�8�=��U�굯���3�yP{��Fөb7T��фne��,zy	[�x_�V����,���Cž�����ag��4��
���E������\}����f����AlQ�S@��B�����=��%`@I�3GC+�Dɚ* T5��a��4�D�� H�%E�V�����%eX'�.؍~2�PiC��՝�zU������'�y������8���b�ru�`z�~N��uP��u���Ο��7U���PV���H�5 n������k��JF�4��iI�z����Du�-�������{�ӽ��kNU����g�Ƭ95��c�ۊxO�Ͻ��ُ4ܧ�%�L��˔�'#@1r~MzXc��h/����&��ft��l0�/2��ur{���66�P�I�h�q!����������w4I�LE�rrb�K+���C��/{^�l��ܳ���7x�+;/�`�~1��9G��;��L��p0������]///���F�+G0�92��n�L��C�'j�K���r��l��rx,ɠ�ig'.���V���ur+��f-����� �߱��^RAe�}��D�E�2mg�?FBt�İ?`��G�f��Ȝ�+��	ܻ�AQz3b��tb�Zة�-�)�����^a@��I����D�`�c�$f��#�.��\w�z{[�',n������ň���L�倿��'k@�F�epF��L��?|l�����J�D/A�X
,�S|(%.A^I�
Ǘ=YX���I
�E�@2��牯�]@luƚ`}�&^��q����-R@m����DDuw�"�Å�*؀�VTV>m�����5�1H�g|ʑ(Z����Tm(W1��O��@���7�t�\[#�2\*j�|�X�T�� 6�%c2�4�=�d�Iخ )��q&�@ 9Ȃ�%����/p|_�8����k;�v���4Z����j8���}��晙���j�[p�#��[���F������A]-���ל� L�ܦP��f�1��j���8ς^�o���T0f=�*�'��wTo���G�(.C6o��m���a|W4�	ɀm���"�/Q2�J��041	�"�\�΢ݱ�c��L�����v�фHe���s���J���r��T��A+�v�٥1�mG��*��P�C��nE����gS�MLL��+]x�����:coR�7�p�����BJ��r�Iti�yX��(�z�֦�4_w#�7�B��6o���'V�����/��q5i��$G)�����8X�X��"��]�o��E��R�+��苡�1gg�Y��� .��B��������W�yP��N���ǜ,1bp�����n��+$Ȅ�j��^�b_��A�Ȩ�K1�
�,W���]���_�?��ȥ���TxiCP�3	5s���jo�N4a`����tR�j������n�o��r�ջG�����WX����ZoD��� G?1�<`�:!fs`˅��}46�t�wt�	�2�����U�J0-{6���9��f�(3��k<����,O�������#���ͱ�5�N�=y�˾b{�w�9�͎�ȝ�=U�C�հ#]$�����Lv����C����1��!.�gT�*�9��t���cJ2�o:(1'ggׁS��o� "zX�e"���w;��&�JJ���Xz��EDj�W���N4Fn�s�#m��P�c�W�4P�Q�V�ܽBbbq�۴_f��W�ڄ���I#M���;C/y�]��3?��8y}}Z���{���l��8�b6�UR,��f��s�s�/7Y��a�$z�����<%%�s1n��_1�l�!��iii3��'H8�*6n���@��a��G8�_�� |�q�lj�+1�����eUlDg%�C<��Z:U���\)e�fgg�{4���|�'��Ϗ�8�8����9�
=����� ��.��c�,\���;O���9|{	�ڃ�~���� g��}Wƨ�� Ui����ss;''��^��|F���P(�+K��@I@;����m�)x俓3��}#Rk*�FՆ��f
LB9ܧ�ু�;�!nf1�}���:�_�;��G�3��uQMNZN���#���"iʭ���B2�	q�8\����+X;��\�H��[�'.�a]gQ�Iaeݸ��@��g5|��1@3���6��c�	��oqc��W���Z0�?H����^���gFL_l Z�U��	�?e�L����t��{��FB ��d?*�\�+�g&M����}����Ȩ�Q~�2I������������9���O��=I&&&�7Tc؈���P0���]y_�~q��t�c 3>-�L;��~�:\/q(DÁ�}�\���+�'Xn"����ݕҥ�/]� W���b�����{�z��*O+r�/:6)H'M��KB��h�\�u{H[M&OA���t�^�0^0��\���qo�ZEpݗ(�Q0R��緕�ݵ�3{|��XO�lDHF.ԍ-+���1��tx�;m�e�D����̽lg��<��B�C�周f���������罰�/Xۤ.���%�' ����;���8�3�Z��2̺eh:4�<���~���	� �`�Ŭ�/ވ��32RO�,"�S{{�Y<2r�>��Z�v ��Y�`���|R��h���~��KM����b�^���y���[�Iн�*��#��Ԛ�܈�+�/@����|����K+%��$tigN�/�sM�N���Ƿ�i�����l��PRr�9�=��)��˾z��eO̡t��ݽ�$Sw�ލ�Y�15�	u�� �77?pr��>�&���W��)_�C��y[U����@	%��h��+y�t͙���5#c�Ml�a�ׄ?�7tMB���E�L�+
�a�ڏs�}7qS���.//�c
N�ʔl������'n���z}�ݠx�%Wd:' ~ȶ��N��ɗ���	Ω?,����&�eБ5,lJ���ۿ��s������T����Ib�u����>��T+~�t��n�Ie��xK,�]y|�OSp��Hb-�M��,����!�͚g�9.T�Ƌ �D��*�J���-f=W�ua�'�oq�ѩ�H���"�+m����*�.�� ��{ו���N�$$%�>��)�X�|����o�ha�_�+�ƽŭ��j`Z��H$*NWK	**��;�c}gOq������/��l%�� ����V��NS3�g���v�\||2�6�a�C�E�~>��d�lAOn�z1G�,]Z������3_�xm�A����Gf�3�K�6�2�f�?D��tRWrIG'�x̉��Q�B��e��?8��0� �a���F�g<�R<[�� ������W��@��HQ�����HI!#J��7�Y���f�2�[�b����AE|��$����JET�ah�W	�ZZ��K���B�Q)�w>�w�p�z^�[c�e54Š���k�δ��*�U�Y�׻M���P�®:m�_���`�ퟲ?H
	E����FR�����Za��x?��)��nT�b�sW_zf�";u֮�������C�s\����t{��(����'AR,�h���_��\�&(\�'��6�X�pÍXF�\�ѣB�W���9:��J=)h�� A:�Y7#�<�4S<�C��q�	��~�ɴۘ���]K�țGT�����
{�� df�~k<�4��uӰz
��^�`���̳���YcG'^�*��N�OK��V��W�;�=�ܺ�=��]��F�����~�AY8v�L�eu�V�t��b�X?������T��j"�텴��$�#� V�KG��W�nk��Od�;`��m9\�n]4�>��E��)���+��Ȅ�E_>��֦���`�R+�ҥ��K���55H���Ygkhj�v�,��`���~��w(�2ɫ�E_���v���G�]�s D�&ܶ�o;���:�N�L4�������������W��$$$[G~��5P�l�鵋/5��21X��(x�E�R=.� �{y�lR<{��F��qf����K��������Y9	���_���pN��61���d}QN�%8���KI\�XU��P�_�������&y6K��z�M�)s*0�x��3Ym��7n|n,��N��;J�$����$.�V [:�����7H�}�U���m��U�"!<4��K-��Ʈ��@{���|��d�⏒R� l�r�Y|�K�r�+~t�o���@��;{@ɼ�O9�����e��Pҝ98`U|W��}Ax��
]�<��z`���Jcm$��t~Y�+-��"�P������������MQ���{,�y��G�����zO�Y�� ;��2 �X���%٘J��Q���`C'�__�uX��++W��wh��W=L{��q��&$S���<���V��I���oQ����C1�W���!��B�8&�7Z�X�dX�Ym1�gm��nք�� ?�+PR�x�:|��3YR�?v��C�]cF��`���-
/)OꉋdNz͟��jԣ(�u��;f��r �9@����ń��_iyU��J�饫k������!9@@,���X���n������vihk�͍�<����ʥ��u:�W �B���A�v�| p�±��E3����������7�U" �}a�� ѫ�����䃓�����+������a��0�%{=%ʛ7��`�/�5T����j���������8v�ŀ���"�M�"��KZ�<��g����Â�>��B�v��	}~�l�\kYѶ�B��}n����?���=޲:�a>��R0�ϟ���Um=��M+��Y�����2�eq���ەy�����ʼ=��Pah��¶��V����}�k��]C�n��8����s{�푝Q8"Q�y�ƾ�g��
['������e�����:���6���mV�苛A$r��:������%��~UD�VL����7��2�˃���|�(~�宀@��a�r�N������Ώ��j�G5����SFG�����|�C��䡀��d����R^Yi���7�y;E�ϸO�m�A��l��V��ss��cRV.�Ý�@���v�����dg�t��\O6!@�A�@M�1�0��_4�b�I���w;�Đ~?��|����)=c���5�^ˇ	�d�����de��釣0�˾R, c�å��q���|��er%�� ��[���5��@9�h���0�E,���B��D`ܾm؎��3J��/���(��ؠL�.v�<�V[~�$���l7�ᗗ7��T��¤���»��λ>��6NK�!!=K�Up2�s�=�J�C2缓@��2%E�C���K���tY��=��ϊl�gGFn	ܻ礮J�Dh�66���\��o|,�L`|Ni���M�3;�--��,����n�� e�d*��,7��Ȟ���w޿� ��4u�����\����x�5��#T !+� �U/
�#H"�����"��S����_.�D^=}%�����i�K����o1���n�,�͗��D 9�ܻ�q�l�:q�OF֧��t$Fs��G��R,�of\$��Sū����c��vKq�i*tb=�y�,
|�L��qXz�EwOD������ݖ�����14M��zv�'	��*G�/�k3�/��˓_�lV�hV��द��n|�ՃV����`��=�BB�Əy�n���Btw��9�E�l�������;����ik��?j$����iȒ�Y;�4��2M�}89qvqu��k���;�mii�GB����$�ܿ�0��[��0`���������]3�_:B̨j�܄X�c�w$UY)��e^h\Q��W�U�V#�^���1|b���B�1����z��8��A��L䘧>�a��qWy(dݚ*�6-,چ�f��/FJ'Uw��#�W�Q�0^��ѭ08l�f7+fW�r����9�g���V)�90�]���g�߈Y�&B�v�{�=�_�=���@iARN��v��d�C�/%�3��!�3�3���3��ȯu��=ր�b��9O_AYY�ڬ+ckd�UU�${���d��NW�x{��|F��CB�*V8~�mI�g���ҠJ���ߊ�c�uDȢۨ�x���?��G	�B���ܟ>}
[Y�I�'�o_Ѯ�=,��ԜxƇ�A`��*�Y�oVU��;s|L|��oJ�&�J�n���[�� %{z�r%�_��4#�����H#��>%��!����"6(��N�~�g#�R����sں'Wg|�7/�j3�	��"��Ӝ�6'�i~�k����Q5�h<��Ƶ���(_�;�R�S�=��n�7-��C�&%�"(G��z:/���`6�!bsp����vCN"K�WIIv��{���T+^P�-��z_��%�ͬ��I\�!wrr2�ћ�����������;�Vܷ�����4��,\]�gV�Rԯ<}:��CM���=�xv%�sV�~Z�����&!��R�Y�D!�g�!ߐ��'i��-^lD_t�n�% Ǘr,1֊��}�Z���29xb]����"�}�h�'���0���^�DR�g���.�$`�|�5
�/C��ҹ\jP�#-1��sƓ������	�C	.�̞��0{X=+��I�w�@V��T�Kr(�ݒV��[u%dEo��j���<*ݡVxT�r�+�\�f�yՀC�^YՌ��z����uq��lZV�� ?�8���}3�?�GnLP�Lk��$b�{ٿ\Z��"U�,�	~��T3��02>�dS[[��X[������
X^�@m �h�s��D]�+���ѥn�u3A�
3_�i*��ttwEF�{�X�=��[��������=@��҇�ݾghMO�"nʸ��C������Wk��B��	Jx���������ʗB�u�K4akDXV�k;o�-���r�@��� ��_V�p�C}���+�4
��hۧx
肍2�a����wb�������o5N�)��{P�s}[<c�խ�81i`�Y.�i��>Vb�W�.���ey.��c��l;ٯ�f�{o[�t�4ɔNm���k������Q �3W�b���+���0UY������'��rSӁ���4�Xʚ���R����FFJ%<�L�D�/�d`�g]b
&O�KF8�>A7� �4��j\��������A����i�XV����ˬ 7q8;^��U��<�]�#Q���]�@I�*��_n�K5@!96����y�	&�Wl�t�Z<-f�]׾�r;U��:.����t��J�*�m��w�uω]�(6"J��QjU%�qo${
�Ԅ�ˍ���?z�J�-X�<8Рk$-t&\��on;B��.k�(����bV6�B���}ڬ�:WW3W�>�UE�;{6Oڂ���/�Q��N���n����;z��k>�0<<�:�h%պ;����pGFCI.("��}���IIX�9���}q.M��<�Ŋ�#b��.����?����J��ޤ[�*Z1Q]�c�M)Zg,ū���J2J���i��G;��mJ"i�#?�j��t��Y���9������)��s\/�n}=�8��ס*'��u�0F�z������0t�ڶ���G�c��ԗ��4�My��Z0a��$�b�xl��ݿ�a�sz-��K3pS�q��0�y���VwOr�c@��b ޠڎ[>S��C�ʎS����nS�323?KE��{V��0�S|:�`8�Խ��OmGo"p&��;�C����16y�L����&�A�'�[�r�I_��l`����5;�+�!
C�6�^�=���--rᕌ.��Qsg� �̪nD+��YS'q�8T�q��q8�89���.���|�n�Rm('���/��\E��hM'u���7���Pj� %[��6e� iWP%��)�� ��ZE��V�5�?,7��U/r��+(�/�+V�ӽ��`a%�$�i��A�\�S��m/��^;h�.(�ԁ����`A���++N���j���΂[�:k�v4�*�������7+�����N�ґR��R�kk$�M �rr^��H?&*{Eܙ�hP�}v�@4+���pI��૥Џ�� �g�x���G�$����rk�,0�ʟ�Kp�Nj|ߣ��yݷ�')\׀�/�<AR�[�@3{o (�PK�M+o�:�P��@Tl<EL(UtA�������ط岏>;r�@��p[����O+�a�M̝��:�v���2�A���EL��b����t�$�k�&?�l�a���Ɂ����g�'�ퟞݿ�
_oS�q�I���V�K6�J�������ihb�9[�t]R���?��3m��'��ܦ��� 	�H(�ʬ�<����N4bo�L�)T�����s!j��KZ�Ǐ�����U�,�uZ'���#& �r�~������A ����zx�3����jb� 0�WK+�g��I$�E��[׊c�@Nלﻌ�c��k�����h o._�g�e7��Ł[Yp����ae����C A��MhI��C�.|"�!���y\j�e?�N�qt�e^m��0�<E�;��������v���.��!�.z9���^��UnS2��U++ī��̀~n�ߚ���؎1�vVK�K;VSu��v3��Ŋ������SF����
)��Z\]j�]S���olr�G=���~ʰsM�i/���P��%z�Κ�L��[R��sD� �ӵ���'&��3y6�߻�V���Z��ߜUmH��MM3o�֑=�6;-�<�C�Aӥ��B~B�=Q�C��Pyդ0�j��֢�#W :A7R?��i����$]Y��Qv�h��Ika{3�OF��rL��'������k2&Kk�)�C�|�޿�32R�1*W@׽c!ë&W��6��W���Û�V���.��B���N�t���c� ���ǂ�穚͛S9�f�\���w���.��|�?�=����<���qu�<姶sj�*T���2Α�T���4�v!./_b�xA�����{KIX��h��D�Y���J	�H��o��b�],Ñ444� *�wi�>pK�^q�cT�O��v�X��A��@��N�hc�}<�vY���ݘx= ��Y��{ ����.���]a��F)���1	�0N�S� D��@�➗v㤡��B�׋�q��Ƶ���x�7m�Y�E�%���&�&���4A����k\ޤ��ש�m�p��Z�u�Zq��oR?�cOp0���>����`zӆ�����/nU�B3A~r�5�i�a㮸V߾�>�Sɝ$s�g��4!}�)��fT1���~�5��; J����Y�M�@l�v���7UG��+a���c�7-���===��9��K;~~�u:��s壗�22��Q� ��_��5�+.�堦�''h~���������f�2L���r ���d�'����>�9���Y<{z�DHx�g|��ѫ7J�z��GG6վ�.�39	�_�`V..�]]][�-v���?
��W���m:>����X��e�N��{0/--E)[�
���l4��0���[���+J:*�����%��@Z�<C3j��H{��=u@�Q��U��+�ŝ��Q/,�<z��m8f-5�����6�RX���=%���o�A��R�n�{{���Đ����6���k��{��~�3I$"��כ*Ƒ�MĐ��#�g��F����A��u�razz���;t����V�Zy�� ���\M�U�|O�$�`x���}a��o22n����Z��~H(�|��&�g/_��^�M�:�h5S�e)�(V�v[6n�*����H��<T������Y&��5��31���k��;S/��Öxl�5p�_ǌ27���(n��J�9S�������%��^�ȽzuR��Ow+��4t�6�Yo�Yqg���"��C{Efzƴw�d��qCU!Ƈ�#���O����D�e�idf�cN%)�Lw�e�է@K��x��O�����<�a�����^�GtmR�>�z^{���4Q8&23憆a#�+H�� �{=������5�7k�[&�<ʳ���pw�M���Qp�v_�l�b�β��i�����Ѓ�\xY���@A�W
^h"��2z��{PTS��DY�?���vݓѳY���Q�m-XV�D�'4�_���������Gf��Hߕm�Ev˱m=N|pq����J���9 ��~������T]9*9����`!s�6]����{��+�]�ٻ�k�t*��Fp�s+(t�jd�h�A�Վ)J05�+�S�9}A]�պv쳾�)�NV�ƃ���3��GȺ7)P�[/��w���q4]�lf� ���K�D�Lc�{��O��UçOm�qqq���$(@8NN�o����}q�~ci�)"%e�����<C~:~�f� ��z[+H��L$����B2���/�N���?���3Ԍ�zzAW��q�,"?��:r¯NO�"�q�v�r�Ɯzff�""#gݛt�F����J�~���Ҍ6�L�[#��Q���.�6	==}GGG�Kr%��K+ ��[u����f�rz�Ҕj��ݔ���M�]Y�����|�yV�XI�B���n��u��u�ؔ��
�>�?���v5Rt=PHJ.��]�,L�9��_��\�+]W�&�O�{�]�����32��I��4Y��/����Ĩ윜���N�^m�/q1ۻ����ѧ�Jf���xSt���y����ۮ��{M>��3ss@��9l?x]9��͍X;O&�iv���v��h:�x*����B��!���#�Yɱ���cdfo�압d{&!�ӡc�8f��]����?y��u�������k���m�Jԧ)����"��yw�<�{�8��k����w�ֲFuR���DH�1T��������R�lT���N����C��f��X�ʾ�j5�,k���2�@�H�M�W�ډ�-d�z��Ӣ�y�g�|��]8��Iĵ;��P�Sa��sqi�Jk�a��]�W��u��JZҋt�9՜�����@VX�$�"�e��E""�&m����h�[�##���34�Ty��	4�y`}M4\H�uE����n��!D�m߾񇇇�㆗�nl0��i6؏P~Q�fl��I�+��,�ֶ�ʦ��#**�{,�=�Z'��ח���W����o������IIt��鮸ջ��θq�Dqё�M�s�����*߻)3Ʊ峩p+~:��	u�����i����ӫB�Sc^�.v�o��B�����t�N%�RYt���+�q��V%=ŠKoP�θ!��<)9S4�=�����	f��.Q�7����;Da\k��<F��9m���k[;�Sn�pYG`p��Ke��,%V�d9�R��z�<����afe�z9=�t$����:�LŮ��(�(b��Q�BaΠh~�26-��n� D3F�oA��hu��F�-���G���?UTl)>��2�@���6p9�Q#f��]�f���_����J\Gj�A������:��ƥ���
��n���xE��Ot����I��h��Z��@����ß
m����*3�'���K��p&u�yh��Y�vfvvB}���%3��8���f�̄X8�>?�^��e/�B�h	T�"�V�p�����dy�������ȗ�Vh�%�m�8��4�2�}�[ƽ��o_U��<��0�Հ�
����+(�a�O#��a�H@O�үyN�&d��u���l>�\'�@��\S5Ӵ�X�fSh�0�sM���2��ۣȾ��������O��^B��㝔i`�������@����Дd�ۢHeKK���M:��_:p����B�f�i�^�����]^P��/)2_:Z8e�7X�GEF�y�p�]$E��R���b1E˔�����宮0ꪢ����Ծ��q�v�]6�©�E�S����_嫪���nlZ�Ԗ��p%Fn~ 0s-�N�?'�ᄜ�Ǵ�!�D��jо�����.|�Lj|mo
���TM�6��k��`l�K�T�M<����̫[Zz��	�#��Xht7��e����.������h���+�&<�ƻ,��0�QvAA��w������v�a=�e��C"��W3M���H��j�{�,[[���"c��wɑ��& �!��Sh��$-7n����ù�1���?B�Fk�C���AoRp����^9�dB3�MOrt��̘��������}�|�٭�͍����Y�/|^�u�.��m�>ZT����QP(���uJ�2�K�HRSD��H�s8���q�@=[��v����!��!��v�*����!�%������V���*�luo �-��*�{�b��GoC���keP�	*	�!~l�1��������k�T��_ut�薹)f�,5L{{yED5��R����%I��dL�G䨓۪���2cC͐-���b�/�М��L=�A�o����}����`��z�TQ�nұ����m��TxhR�DP_b�ld��yH�f�)tp��>���E#ߍ��ǌ�pӥ孺D����	���}�c٪�5i������5�K.�rbi���S.�(	��)��ʏ��i���3j_dӵtg����A�+���5+/g��XR����9�Eu�v�H��`� �&�"eÜ���2ܟ"		y���C�UL�<h|��.��5�ς�p�8��%��Eb��]]���yGvk�������W65E��Z��@C��x�uXՌ絘��J��Ķ�k:H�����WJp���d���o
�N)��wG�A�:0Ӕ�q	�k�<oE�8�PS�n�Ȃ� =��^�c:a5F�o�����IRdZ{Kg�!���l�ۋ�w�*��T�<b}u��@�cx�ו������e`,�h"i�	a`�;(��J�:���jE��$����n�<�n(..�QgN�^��_�qKU_TNNď�ؑ����XJGw�D�=��s�	k��q)�������n���F��9>(Ywq�����KK�����v�=���O,w��ma���&($��Pཐ*��t�D�ľ+�8V�oZ���n�ݓ^]��y��q�8B��C���ʶ�ë1�J���@��W�w{�(��|�^�+si��C1����q����\�ӥл�Vj\
��-l�׾>���̸���5�%�G��?��h�Ԏ���5O��4o�(��:	�N2�\N{�A��G�-v��.�ywy��P *I�����L�����+M�U��my������������:Vu��K����D�#�iO��R$�g|�$Pi'��M��63<<#��Ɠ�0	�<~^��?E8Y�<w��2�~t�bP̃:�j��o��>]�@/����~��S�N��P���J�k�)xv���z�>?��.�\c��O��"�����gΠ���
�#��P�N�������&�4�ʉ�B�?���93��a�]�%�u
ݦ�-���χF��ǵ�c��qо�+�Zwň������Ԑa4��O�@lԍ���Q*����y4��_x��Э�;=���׾Z���A!*)���}*@ղ�\L������b�(ik�/����7=mű�S��T@HDTU��X:0�Dx}����9��l���^��J�>����� )�L�+Ƿ�:wr�����Ӄݵ�،��&ip�M�Y�$%��z�1)ƥ ǵ��������3�������;��շ=�Z�w��oy�=HS�V�ֻ�d!%��0���c%��\�R��7X����b�͞.i���)td�P�n_�����@���N�9�C%L��6aj�3P��
q�9��T�����
y��~���>�+��<>Й���p���ϘO�Q�XZwvb��ʝM>T+�fP�߿o�D䙧!Cڠ~��=-��n�y�r�O��.2�� C�*�ƜN7Goo��ǅ=�#�ӣ�����I����k2U�b_eJEF�t�����3SVM8u��;hX�I>�]|�=!B��A.�%-#!a|QRr����_�
"`.!��zt����Ǻf���?�1�y�(�9��^�(>����N�f�d�K�+)���-����ND��:0�
|,wo]��g�~r[���,� �}��h8�p�Jf��Q�-���+WWe�ˠ�A�vL�զ��,�J�u��� ��}�wո���*w���?>��=h����5!�By%H���{�%3��������OdZ"��D G�-BH�-�i[cFM��V��hȡ�;8 �'wF?'ٽ�,h_t�D�,IV=#���;�^H�B�����zs�b�I�3Ow� dE��3��kj)v��0�Z#8�P<Է@�X�XIPq$��R��Ή�8�sR�}�k�c*�6�����ts�"��+�'CyZ�t�t��(X��E���{��ɠ�U턜����ǵs1j��]����nn�S_	�G�g񀘥m�=#--lp��|��Y�n��(�6�=�-�,��xH�ع���T;ji+�u���� -\\��	������TH9:�	[�D &  ���N(h�?�42�{B|9�.JJ�_f3D�4;c)9W���wr�e�y�Z�Y���|򭎯���U#@Xٞ�w�a��z�)��2��V9�F�CfC�#1�����Z�G���g#mH44�����/����g��~ީ���f��������|Fژ������\��"p:�[������K��N{�`��f��@���}���|�[���I��/N&�P;|k�r���,�\��9�b��	���b�7W��;������Ā��w>�j�!? �.�gܨ��G>�b4��㡆��e�s�WRh�|�zն?�MZp�R$a�_��6U��{#kG>�ZvH$Yt�X��p���0A���/#5>��s��<��C�x����}8���p�������Ǹ�r�UH�RL�`��`�@N��3�����^Q
mJ���k*����g�[�Hķ�A@��ܑ��.z��|	��<{.�055��	���{\U�q�n?sb��Y�p��t�0>|��<�� ��dG���S�Y��
1��T�֛�6���jrh�۲��4ҧT�9w�'����;�*Dޢ������L�$��ȸ�$�kp��S!ޓ��5f��x�cr-u%~:����@�@�Ix�@M�\�u�2ի@�o�z��ғQRާ�uK�����Yg./�e+��%M˸�Cw䋮����)4��ʛ��S�l��gTԽ��١�ˀ��/��DLWpZ������ϘؠbX!а�� 4���C	�̞���`T����^Z���qq��L���ꠅ������?�Ro�Z��$z<g���I�9Z�G���4:\�b�
t)Q����"�3��=�������̖w�I��X��> �K�|��E8~���?F	������yJdh;��
_�������^�����fN��O#��{ ��������W_:����n���E��x�>���ˠ�{��MV��I+^-�J��m�6Z��<M��ށ�k�|�2��"����N��ڰ:�#l:�<Iz9x�[VI_x����u�7�o�bt,ʥ�ߠP7}���JJ�:�1HNFv2Z߄��K��������)�%%�15�y^6��^0ۗ�r�W{~��u�O�ࣖͰ�C�F@@>� U���l�gd̅M(Zk'NA8x�,���+�Ag+���RR�5R8�&�Fȓ�LFQ����i �Ϋ,rd�O'�?4wݗ��휡wʎ�����o��g<�G���I�Aֶ�AV�ʉ�@Ĉ��B�d����M��>�:����k3��I6Y��H-o�9�=Ar8��[[<)��8p�������x{�֗���&_���TR����D\A��ý�ۀ߻�x;��w�:���_Y�"Ѐ��)죦�(͢"���&���dH��
�4'Y�Fn4�'%=&���L�w�SU���zxuk��RU��A��7�_�(�1D�0%G�%V��4���
�:/�&R�`�7T�|Ñ/ܙ�l�����Z"��=�H�P�C����PS���ʅ̂�@l�u�l'�F�?����Ύ��;WMm�~����7�V䑙(�������f�,ll���A�
�M��KemoO�S�����3F���e�E��7��2���g��k�c�SH*b���k�dq�p�AS�C�DC��A���|_�6E ږ�{khh�$KJfA������嫠�=:�딀���������P�J>#4��2��v?��RzҤ�$Ǭ��%���!��R��A����a�1�q)���#����*#�B~�1�O%Y�/���}W���z>���Qndf��lBl�=�c�0aɌ~�3ʋd�+��Vp	|�d��1�E��EQ�#����ݑ̐�������g���`�"�d\������{.,�(�Ʀ���!�΄�9��'�@�����f)}�;M|!�ijn���ε�y�bi)İ�5G�wvB��YOt5*�լ,�������2�cE*�yt)��D�_���;�� [�����r܉<z����-H/4C������=�ݨ�r�ڹ��%O$��;фߘ�j�Q6��:p�|�(mB��tyX�[Ф���_�@x���X��_U��vw�`R�m�����0_�4�5i(�£�����?��`�j��ꭙޤ{��,ͧ��˹Is!j���m�|8��n3�Iw��}ĺھ<���O��śĬ�Ak�x#��ۮ�e�9p���v�+:S�\� ��f)Z=~�\3>���/����WKK�����鞒1�3�y�s);�G�uu�S��k(�b��W �ݾ��r*gPl����en[e*�x��>�T����uM��HuUCK,S���;8s��x�wq�!;p�u�%,�"�@��/�ފ������� 6^�dMB#힘&Ĳ7���}�������NJ���P�!�?�}�t3�w�y��Ś�?�fe-�~�al�j;d��v/f�	��i���2�C�P�����kFFС������p������g��0�(�|�@tpb���f�3��n����(��(P��E�D<ˮ�P�9�{G��`��w�''a�koݴ�? '��G"wTe�u$�߸
�ii���G�y<3o�%�K���HNLIq^(w�r;��I��#�d~�
��׻�LӲﴙu�N������K����7O��4�)��}T��� �Ȕy��
��-j�A���!bCF7��no�nz�ה�`�X^Ǯ�Ft��\�Q�Z�?V���Gll�ۓA�EH����X(i&%���WcV����b����;�8Bŀ��F� ���hfU�m��/6�li�C0&�QG�Ë���(()Ü�Tg�]&�`!�� ��$ ��J�(���,L��n�2IN %�O�rp�M�F��@=6�.�=ͳ�[\��x����d�\n.*��(:g�_�!�M[,Mh���$�>�?���0�D����L:S�������@�a���-b<.~=�pff����1qzA�>~��Θ����c)�	+,v���t����~ĸ�q�SS�C��/(�eQ�Aw��	��Բ�g�y|�Y�d��=��[8��u}���97��>k1WPXh]喾���M>%o�J���㒕�M�Ѱ��C*����	�+1�y��H}��kd��o+�"�"6�җ�m�&�|Gp�mk�2k?x���y��������j����:�&MM�zHr!4
�©�e�>fP<��>7���k�;��iďZ�-(|BE������O��A�.���es{���a��_�U_�FSrLnYߠb/1.5�8���6����v�?Њ���aVt'g���
�.��Uo�z��Xw�Iev�RU�����}B3B�����a�be�* k�i�§=�
��v���B�����5UvD�I��.@��u�Ɯ�_���W���w4E���US]v��+t����ܿ�}��A�mȰ�En��Puu���I|�������A����w������GC�H,����rPKqD�0f��bb�芖TϢ#�Y-�\ǔ����o�B�����k��ލ��O���_&�B9j|�+rm�#ǋ�B�M�feл�|(����6�כ��>�Xp���P���\\s��U���)�n����3@6��A	�.�Rj$��6�EI����Z�rn�|a�����A#RN`$n�N��5t�l�m���7X�TE�ƺo�zV����C��&N�h^�Frh�*����樽�G��32X��O"����o������iۉ���r�;�<��J�h!:��u,�MLxI�����wd�����[cu�^��W8��z)Y����Er��=�T.�et@Gm?tG�!�\8fd��rÓ�kHj�-_Q(�G`{�a���7��  ��}�'<��Pp�O��S���^���4�N��� ��5.�����\\o*��Z��������e:�����W�R�����Ç�;�z�w㔄-~�����i���~v;��ú����C�ml�S��F��2q�f�b����HScy���z��]���Ϊ��r��jnO�P�|�YD9�$!$�>>.�םb�C�V}�Z����"��+"%Ek+�B,q��^�^^�qj��n��G��bT����Մ#�C�����G`��s��(od�C&Q#��~��~��� T�k��jb�&H��:��#"�kv5x8���J3ā��fmӔ�J��ZJ�T��~	)G��b�w������������o֣߮�z�w7�e+�~���8�5`�|��\��
����j�h�0��B]�����}z�w�L hZ91�yLI�C����c��b��g����[�u5�[�������<Y��� ד�1�
��LDD4l�<x���}�4`c�l����-N>�����I���'�踴��-s<},��?��r�L~�X��]�]�U�T�8�v�;o�J�*�Ƭ��x����l��e���=�������.7��"�ւZ��j�i�[" .c}��-<f��[&ER�W�H4]W(�.���:�r�����3XT-4�tlE�.�M	��n��ncن�5O��޺իF� ��iZ�Ĺ������ݿ�Ƀ�(��͝�ۿ��#>$|1�^nF]*�k`�ƋXR���y��b�j̔���[�z�|��Q�Yx��;-^P����݇�'�^�Q�����]pR�?��߷n��i��W�������=�r����ǜ���A�{$��Y�6�p�-'U)�\����|��Nt�b2���[���Z[K������
�¢�}i�wJ�W�t��N�a�� ��H�d�Ι����ˋM�L��]8�T��֞��w�V���_κ`Fƻi�)�Z��+C̕��ۀ0��d��!��-.~�p�Q/�gmv�nG��V�IB���&�,��HYA:�uٻ��O���?��ʏ�md��\&H�ƜN)���6j��u���mo�0,���E">ߣ�"-��AG�1�F�fcnF��K������z� u�4-^-�AR��Cy�N��^o [11�q���b?�S=4�<`��e�����_�3t�:W*wn�'���g�R˰ B�Ѣ�/�%?	����B����7�}tG]\�>;<�_�|������:5�y�H_;�. ���"eGX!x6���ȕ*"�u%�	����@Ha\��8��]:3U@w�G��o�z�|+���9֥"�u$	�]~�ʝ�V��w�!�67#7}J�:1�A�L��"W_
��=ٔ�7�{�\�9�'`?��!4���z��t��?_Ҷ���iQqP	@�ٙ�C	�=�fzI��.��B��<�L��[��R���T`�w���(���xRcVU��f\z�z���T�����n��\?]c�S+�sH)�ܰ����Tb�)W_��g����q.A��W.��0.�]qI�E�b懲�u(F��ȗ�CM7��wPr}u����e��G V�)5�}8�����!U ��LLL R�f?q~���=s]?V"��,q��QE�$�O�ax�K�=<҈Jau�� `��p��טG�G�v��z�;Y'k�?C
HjŎl�D�IE3nŋg�6;����=��SH3h-�A�Mդ��%BSU>Ħj�?�0i(���#٫���z�%L����3^
zƿx�IU�I����1�Rv�oA+�)�CZAs�zA�n��6��Ӹk-71s��QiJ9̂z��knV��;T��c��qmU�(�KJJ
+l>G�@g�|����{ﹰDs�+��{\a�o��� �#�@;�T6�\-3��>,n1b�����i�; ��JM� �á#):��e�ML~:y�g���i��
�5f��^��)w6E ��:6/D:u��uȻмoc9)aq7a~N�XY����)�WS�9N���5�2bc#�Ԇ��5A�)?�kG���m�t�e;�θ����d�!��(���s�:���'F1��:x����zo�]6�8�3"MGW��#`3��F]������7�$/������eƤ�e Es�����edd�Û���g�G�G�����''lϦ�"�oo t���!8�"K��b�H�y��T��IPP��P�I�w�.��	��h��ѱ�/�Ņ�+��=;ğ �,x~�C�@5���䤗R����8Pz�S��[���E.�RѴ�������s����ɂ�[U^]����gV�=�!������^o�˟#>'v �{�4��))(>��(G-	⭪z�ܰ�v����n��	7�9Jw7�f���o�9V~'W-��F���*�<uy����!-�+-��c���Gm��+)$���Y�l�V�w��v}���gc]�yA������{{�u>�ƈ��<��:*ѫ�#�J[�������"��DЖ'j��e�+��v�mjw��cɉP��	.4ꥸ��pVK�b<�U'b��S
�P��?;o�k'���OACy�� �Ӫ�o���"�lR~=�~hXj��N!i��a]�q��<t5W?hߏIp�gc�}����*eoo?��؜��Ԯ3��!����wHbk;g���2��5����Ejdd�X��F�c���+�-��Ⱪ"� ,v������� �g��tt��Ș_G7�Ck��qn!��)Q~z���Zn�g�9�ɖ���"s��&�*�?47�Z���{v��9,��X�*�WJV��PR�Vq4�E94�9՜�6�{5&��n_�3��~�LO}Z��O\:���{�g�`�C����P�����6��ه|al3�?�^������I������3�;�)�(()_k^C�4�
��*_��OL<���%·r��=�"	D���#Vټ5O��ʘW�ZW�X	`fUU�P�&4K���i�%�E��S�0��s�P�0��:|�L�KK1�9�L,,��by&Tj1.ė��"�d�/�dx)�/�5`�O�/��w�/F
�C�q�_�|��]�u��]H��DT�;xQ`P��T�%��֭4-��Pg�|�0R�2�#:�%��Ӵ�!���I��@�P�,�<9� ������*�O`����b_'�E�b�v�׳��A���k��px��Wcb��d�#��lWUF�6���������>���t�aZ���@A*#�3�}7t��j@)�)��'i�XIz>S3y������1|9�F������� �Jfx��|	D�����*_�>:���h!�j�ܜ������H_�]��;	hq#?o���j��U�N��ʙ���^~�����m�}���E��^����m�
��*�q|���'�����!�&�4����Ҩ�K@��D��ԄԶ�V��.a.��А�4�&]YY��� �A�����z�/	y�K	=�w�B`\8o8*ιIS�TŠ��h9��I�b`r

���!ó@0��rCS��n�9�[ނ���[��B����wO{DV�f��q�]�5DZ�mO��������?KY�	y}��#�r�p���z�mH �����ԤW��VGˀm��8U�s43颰{�K�<���%Yu2%�6+�)�}�FKt��d4|-S����y�����o����^TZt'�$	�R�R��~����^���INj�,W��I:�k��������J��9www�t��[\�1��I�w���\޴�����
AK�5���΀G%�K��|�]j���'c�܉�׫9�4��1~�2�?�91'/n]�|��ɍ͓�c�"��~�iB�Z*|pMsꚟOFbgf���ř��Hl����ǜ@�zhF�|��O�����~I��]�g��x�|`p��]|d$�ڦ*��2��ݫ��@a&�Z��y�;��a��KF�j===�H�9��"��T���'dn[;A��G��Sw=iVx�""$.ŧ��G�6�q�{� �ԩ����JB��7�*ӳ��z@*|i���7�O���p�E-M\
�[��p����������U�5����_ye��VH��[X{�J����oət����\��\̠J��~���4��Ԥz���t\���Z�T�5Q��`E�\9�I�B�+��)��Pq���
��	�B�y��k����&8���'��_��߿�A�W07��eb��/7��e��R��1�DR^F�Z��Kr����/����i?��5�ξR?�"���P52��?�-���p�����!K�9����|��cH�6�
G��pr�'i��Q-�����s���݄uP��=���������J�*�O����55A1�0�����-Z�(�*pЂ�F�}>�b/7בmaa!^�}�s[�P�R󽳲���1�.UO��m��Gf<pB99I��x�4Q���� ���̀�u9�h'��Q�^��_�NiX"3:�����R겙)�޹R�l,w��/]^4��u��(��Y��i&>�ٱ���T��+�
�=���n���_���u��-��ݣ<"r�:������DԤ��qR��G��ח�f���ۖ��A�"��$b��������C�Q��{�0��r�aQ�����.�^�������M���%�[�hh�ɠH;��UMMןS_�"	#ׄ�.(4���75��Y�7(�צ-gfa�n�w_�}F���
��o����Jv/.���BU?�tZ�`��SDCM�p	�J��#�?��wB�w���L
�<|IuKU�re�枸��8�Gd�ڽ	xR�,�BY&4����Gh���7|��'���z����Y��C;'� �	h�+ ���J�=,���>=vL
���I�h����Es|����axw^�Ź�KEh ��&��""�X���(Ɋ��hi+,L��x>�5+��15�:�H��4���̴eZ�(�K%Իܡ���v{qw ��(���%����xH8}Rx~��b�w$[=���cڹ��8��x���u��e:-29�	�O�D�`.��Gr�F�<���C����v	�a>�ԏ8�ډ[�����m�0�\,q��)w?��Y=}J�P��:ڧ׵��q���Ʊɘ�Ɣe�aj�Dj��-���v�����^���t��%c����2˲-SSc���R�V�R�/q�{{1:#&FR���.���Ѥ�{ۦꝲ#,D��3w�Ծ��§�/��aM��^�鬟K�
�`h!��b��O�́���+�3���C˪9[��s8if��j�f�[�I�^�$��F���NN�ߪ�{`�o������ʱq q�J���{�eDR6.&�Q9J��M`[n0.[Xx\���_>�wH��M�&D�_��7�,��^GF~Ө_PzX;����S���eR"5�st$ ��\[Zbj���/�Ё�v��B+�C�KJ�e���mk�n�˻�������Qq\�_-�k⚰�?&���5i�|.Vd�5c]�=^�P����)�J��?��Kّ��?�r\�d�2��!���κqG��v������w@N����F�©�?��d�Ƭ�N��X���N�Q��a��}x��a=�b����3�G8� $�Z��{���,��o�+�d�jM41]U_���6E8B���X(h���
!�����;��jtu-2��d۷�\.(��Pc6\32r[�]3�H���b]hi�!M\�����&�����y��e8'�W���[�j���Q�6]��Vdƃ�a,�4-�����E�t����Z1�>mr9��Z`|�W��Z=���6��a�ݽ�Vʹ�v�c
^JfXS�Q��G�jk'����'���������k�	!�m�z�G����|�����K4G���@@�-�gfޤ��-�<�Icg��.u�پ:H7KqSJ����	l�ņSS? ��'��y�Ȗ1�ħ�
M���Q�,��AZ�w*Ãc�!.������1W::�	��4�[�ir���5�u�NsH�҆��e�)��߳󭕪ܚN��Q�w&r�=�)���Ż�S.��g3�RvR��7�W����UMlC��R�a	_�޹ YcN��<�:�>>��
����Y�|�I����c��{���C��/��r��l��){�n�������JJ�s@���=�i,���!����wh�WU1pr�yvK�b�l͞(�b4c�9�m,A)񇠤�Sb���=:�����L��_�aۆ���!mxl��Q�,�ٟo�ko7дC�)u��q�uSoD_�\��A�����L�Z��K�G��Ӥ�3��͞8i�{mp�3��!���.����i�FC�߭���GЛ����	SP-̾NL��`�Y[�����S�%γ�i,�P�BLX�Ga�E,�g��<a�;Q��Kz7j�n
����v&�5��>���'r�Jڏ4d�G��;+���������;��Y�0�ͅ�l��.e�� �S4�_��ABs����=�C�$G��j�R��c]��mn��"Ɖ��?ؒ�1k�s���dT�҇��AXFW�w\jU�� �=ʼ.�B�!���)v�3O�wS�R	���4u���!���~�H���F�;�/�-�fҁz:�l�$��eirg�_ɺ�0�黹��E"�1�++�"o�^6)6���q�2�Ihw��K�Z6�o
\��Ov__��Gk>�oA��TP�����q|�"�t9��֖��i^���d�d �
�9?CNFF�ɂ����yf�5�Y2���v�-����
��Qp��%��]���=%K���<$P��"��mP'�}� o[�2'כ�Q<lJ��@�k+�c#U��Q����}����S[��.�9�韭G�B����dZ���{]E{ ƭc]M���2�1����Ɯ){+��$�p��Υ�]sK�g�>M�|��b7�r�Z{6�����,��ޕj�+k0{&�HT�%nS��[dbh�����{5�ܾ]H�|� Hc�		�΀�G
G  R�@�x�3	��o<P��Ⱥ[$�,�A�km�"�8�=�����u
�F��+�f>O�f��_�Τ+Z�E���qY����Z,�mjty�**��2�Xo��o �$i��V�q��4���ͅC����i�#v��@d������M���sjc<��m�TP M�r�2���W}~s�ב>�..l�^�H���nj�$$Q�GT(��,���Q���'�޽[}.��B���r@y�MP�������֡q)�Ck��ԋ߿>�x�s�/�@^������;|����Z�e�~���%���f���tk��i.�z�#�y��g�ܿ��{N�e��*�Y2p$�Q'uom?�lè�h9��l�yDV�v��?-P�W0�o�y�=�g�k�YY��a\�Ω�{T'a��k۷�f��k��������p;�����;��;��7B0�C?ڣy�f^�"\@6P%���<s�)��h�Jp0Ć-��ؙK�l|JI1�[q�QW�x;z����>����a0R���-�~G:��gci�©]h�������� �X82uX���%tt��ϥ�o��7�6�g+nR	0�N��MV���NM�rr�f���2uH���~��w|�4���,h}_l���q��qZU����Cp��U����:~'���yOu��'�qq����y���BxJ�J�
?�XwB�?���]O*֏���ww�"|��3�V$��c��a�Jk1�A�����E������9�G]�]GǇ�jh�g�������$G_~1.�~��y�~�R&SD��m����ƀS's�6�jZ#�a��^�"7�h���a�P=�D�ӛ��??D�϶+�SL�{���d�F��<�o�ڱT��ToI��@3u
sͫ+�N䮑�f��,�Mcޝ��u��C�|��\Q���D����x���� b�f:�RO摢���3/�����ǎ���� Y5uO�Cި�g���c�����j����WUz�ȿ���|�����=z�(� �=[n��i�{�9x���߆\k��-H���r&�*S�ۏ&YL�<Q ��g�@2��`n@��:��fk[�:�xo�[�� �2�@D	�v��DY5�3 � �[b���h\4⏿"�H�Oh�
��V�S��(��σ@u.�8R�E6W�#��lE���Z�<�ԕ6^L�&��[9�zPS]���ƺ�\��)�ᑾ�7�߿ �{>���s��(!5�BjiϠ8�iVAABq��"x.9����n�a�[^î�Ы���\����N�����_"�O�C��$�F����%�myNz�70���J�a���������m<`�'KꖜL�{���r'�fwq�K��=�SIA
�~�5��u%>~4�7;ED�=#qhA�l�G���2Vf�����yP�ŉT~�ٛ��ba�"/¸|~�x�27���������i*)�6ݻpx�_Dd��ߎ;�WZS�H�LEI
 �@u_������*��2z�J��������	zu������Y&��C����L����E,�^��Ϧc���h/t6kd��ODD�r���(�f.�?~֠iĐSM��Q���hypȽ���,i%V��-���E��B�O������?z��J42.���j���i�x��@]>��h[^�r�����Z�q�1���18��0�ԮZfA&��Q���1)eX���*��G��d�UWjN��1'�yv�RW�ć`q���iI�CK�m�|+�X���
4 !vf8-�����m$j��)�f��-Ⱦ>T��}���Q)��[B8_J��4�qy��{�[6@�p8�l�{}���@�uzZZ[cVۚ'��%��֘��̿�����k����CH8ۋ��Z����73o� ]���6��Hj)����Xeq����~N���q�K�<��QFbAE�{�����M.��O>���W���혤����9�A�-x���A�O��$�#X��=�V��;zs8����h������g_�:�)��J��E�yU��<+��e���"_3ss)WJh�M�"����y�!3�%��aSo�
�.�`�{}ccg�T�*]��ڄ%�#;੟H�bG���nK���:1�|�o�3�*�Y�#�|�	���j*�55Qj��徛�A3�2v�Z�q���J�<$�,��Z��ӳĜ�$�:�K��ۇ�Kfeo��W�Pu��1��7K\���d�9��߹���ڗM����������J�:��O���N\�d|����Yk����UP�z^!�F�lsII�L�97�N���֏Q�u�.2&;��ɒ���}�N�8yc!�\��O]���%d��q8{ߏ��K0� ��Ͷ6��&�>�����W76�_�/vw+|�x�Μ��A�DW_�H�ΨN!iG�z�9
51����Qg.LZ���������˱tM�G��J�[8~j��N�*S�}�<��≵�!�؆�*F��u���x��	D�2�B#�������^2��]���h����?7ܤ�-I�8/�{D<�4�������^��F��%p��x͈{;����[|��	?M��T�����v+��������=����P�L���oxXl}*�E-·��Ts7��0(�)?y���t��rr~�c���&��3�]\�i�aw�}*/O���7N&��_�� ��X��jl��3U������d�v�a�g��������c��rܷ���%��h����bB�I}�>�0y��r��!s�/��WnG>G����|��x�G�?y�h��Z�}uHH/���������~7��{�M���kb+ѻD�ND�-D����G��-�[�&�FD�D�[��}�s�8�e<c<�^�Zs^�k��ֺM��$W�PM[���������[g4 ������kt�6�9�����cOψ�h�h�\��@'�)tR�X�if�7X2,N�+p�c��� Y^C��Wޓ��i�^)H�[Ě��	x���ѡ��(9��(�7�74pm�\���n�R�$�~������Iz�|���_�����X:
!qJ�J��,֏��2V����Pm̘k۸!f�Y���̾��!��I�L W�Ұ�S��b��I�Ќ���dM��{�:=������`�k�X�Ew,';�Qx��
��@��W�KH`��D#�d;��#L��C�Q��s;�󬽋��gZ�z�3n�8�3I�;�1;�mW>?��R�^��$�"i��pK���t��QSW����J�����q"�6+*<Z'l��`e���0���q���\��ҙ�T���G&�(ǒ[RUђ(�Ճ&ߔX��U�� -��iN�\ނ���S��b�੼`��SD�c�*"G��R�c�T�h�ݦד�ԒI&~����nlz�y���G�t���h�xң���*ݘǔb���tGg]�������#����o�v��7ˡsT�e�sM+ӌ�����ҧa��{w�'�N�bï�I6���i1��c���/�F��N~=���Kx8�?A�T �����l�������ߗ�`�+�~����;���[y�+���g��"ECz2��/��������)1�SY䐺�o~��O�}��פ�xd�z�������=̽9~����A����:��ݝ���L.o�9i�O�vk�u.�8�xB��1�R��8@���ˌ[M�J?W%:�6@7�MM��*/��:�5�7�-Gj��9({s;�'����݄;֙������M��4�i�i+�hiU���-���X�'IQ3j�HQ�i�c���:�[c/���7� Ij�c���L+0�ؐ.�0v��T3��]x������s�Qӓ����^+�Sh��s6gf�Dn�N���,�]xe�Dal<�rtûYLra�� ���K�}��`x��<�����gP��F�jλ�m�{��AKX���P�{Ѧ�
��GV0i.m���Ğm4��6��f5 s��Zl���][�O����8����ո����� 
7�;:�:��s�tv�y��of��uv�*�Sz7.�#�:C�,�u.�<oSsQE��� ����LK6GD,K�ᐓ��:�;��R6g����\����5�z�.�/�~^9mv}ƙ��ӥ�T�@����t���Cf�A�â�����6*[���mEYs󏉷oΆ����}�l6���K��5�]k�O]b�?{����oZ�q�2p�	������T��h���'�j�v^�O��2xJd���@����47�U<~2i~�C���F�lU��J��Q{�VI�u~�FSk��t�t�uG�=)�����d��X�O3H:�݄�/Da�
���� R�D5��8Gt�H�Я���\9����-��L�L����;��}!��  sQ�oJ��=up���%��2�����w� ���T�؊ê�v;��9��~��������2���=����h�`���)Ѐ��k�vt\|<Q9ɫ�;/X�xn��xkr7�G��w�I3yJ�N	K�n�
N(L��q4OM���Sl���Č��[D��� �CN�!~fi��֚4ɞ����A�AΛ�Ɗ2���c��K<�
�XJ("��v�g�t�i�f�7c4y��$U�{�/fc�S��#T�W� �g�=֋m�10pG2��_ں���NM�$���%���D�n�w4�8������QJ��ȵ�c���B��|4PȷX�|�& ԡ� #���3�9u�����?Db��_��~&� �r���I*Y�ʊ��9W#���E��n���S�Rn'��N�k�f�����P��v������$_�W�D/���0�8[�x���c5�59�Td��Ԇ��anT�v����?���ha��s�zn,z��D��x��S(ӋFP����jUlf�|�###�����>Ûvu���y�v��ؚi�-�h*?���*fi>7�V��m8����a���;�[�%bP�Ҹ��W__�R �8���p����$�}#������*�4UD�L��`Y� �B�s��M�"����[�q�KȰ��As��bX��N�EG����K�Y(p?�����۲�ɂR)�, ;"���T|D�]�?Bp�V��U�EI	7�����?�@������/��ݓ��񕑕%̶x��񫑒vY))�� m���yx�vɓ��z��쑹�t���M )�]���/fFFK��R��I�����F|��E���~s�aċP�b��~EZjꗓ��
�����=���]�)g�o�ɉ	n	F/|�r� z���o+[gm���1M�cR�׼���w�&����F�}c��!���{��+,b���e��hN�ui�B!G����F�Cz�<�C�J@��D�2��>(����h����$'�Dm@�paa�=Y�Jc�	r�O	―~����1p��C��b0KVỈw��y^��������m�[�����Q�S�o��_]�Q`5�I��r6�:�ƗL���M��3�CJ�W$������?�r��1�G�<%��lu�q榕������sˮ&!��s� ���h ��ö�N0)_�$e}5h�G��dN���X;n>.p���]����41���׵��CJ�vE���///O���q�& ��Z4�a�n0����~�@@�����G;�=]�;�>i�B� �s�������N��_NL�Ȱ��P|�*G�o���*-�x'CF^&�-������f�b����/�bwd�wvh�<2��-��rۿ�Zߊ83H0���<�9�`��0���І�~=��wvt�֗N�s�$��Ls;l1�7|������#�T{X��5�ʓ��i6�D�H���5	�M��ޅ�����`��KX�jq�u@�+���P�O6$%(i:��n	8|����ǜ+f�v�u׆�䤘����nm�n���z�#���~����
��+n����䎊�''��ι�{y�F���9�&�]X�v�W
�0 ?b�(�
���`A�W#Uo3*�ڪ:�DSK4�J{&�sx������wu���k$��ro��h��w��z���	H��:�ߗz,�� �$6��H<�>ʴ����r��!&�Ud�%���Q0�oo��آZPa���C�1�`r򉘌��-�p�q���l���ߗE~o�|�<�Ё4ޣݗRCSs�I$���o�|�3��V�XV�wK�4�j(e���u���H&��Y�n��}7퐊�.�R�#�}c�v^!:�8}����8�&�e4Ի�o�m�U��B��-T�"Uoc��(�LIM}�N�]a��[*���fff���)
p�nˑ��I*
R�s#��$LR/
K�_��,�� ����� �)�c�QC#N�"
,��"�S]s�3����Xݒ�nnx̴_�'_D-K�����ˌ��2?�6*�?k�h,$*:W���߽0`�C�mF����G�9�]�pg��A���۫������j�G�s��B��Nea��r��%��M��D>޷
t�FmH�c�ٱ�{ˌ� ���T�v���У����cct �������L[s����s�Ƅ��yU�{&�]|]
�]�����@�K8��1\�oW�`.��������lL�b�W��g�M�
��hL>c#G�r��{'�JJ��h���7u=�o�\��x�,���/XD����=�#��˳&���M7*ߥXMx�HC�"�g�T��ERcF����|���w���T���U��夘e*���R��a��C��]ϦnB�	'�y�4�_Ic���K�x�4b�/95�'w�-ڀmLΑ����&1X�j`�#>���ޜ~�ez�K}��%�B�b��ȵ��(��^�(�_�'�ݹS��������B��`T:@{	�g��Z�0R�im�C��sg
��c������` ���@����#O���m�(.(����|�nEz��*�6f�/�v�~��~���������M�Q�����KV�;+*�x20�?�&0��Iʗ=X�n�j�罯��,���Ƌ��1՘R)�ć��>��ݳR"溔��(���R�O4>��2�Kd��~c��a#�fUX͊�?'�ޡ9܁daN��r2a��4���C�� �{ﮩ}.���v�9~G���?�;"�+-�S�C�Qp��,��C����o��k(2��ܸ��}�]x������cMr�?��l�G�?VZl0��ueD]S��\��e�փ�P���W�O;/5Wd#����7..��IH��eE����>�ԕ��nN7��+x>�|�{|o����h�ܵ���w�ܡֳtY٧k��s8;{�W��H��԰"�r�{��+1�B<D"Fi�?�*�:z{���m�}�-|0բ��ՑZW�\�%�m\&�ø
D*�4��kN����G��i�=�f-�:5�$ҳS�S���y/�B�9���c) |�bꂕw��/߿���8�:
��XQ�\V��MHȓ{`�������S�����ݫ����C+)���&t���u/���M�UKo�Ͽ�����(��~l�ٮz7�n�����ѳ�f;&{�+Ū���9�(�okk�5�1���VEߋ�^���z7�Y�8[���3��140j�G4d	P��^��w��XG������S5�����EҨ�1�$_cF�d����?Ժ6���{�Ux7|å��^�5`����X����[�ty�4��݄���_Ye����J�.?���,z��h m%����%1qq2�t;��¢9�]��55���"��b�?~�4�6$�b�^�����rQ�~_~#3)A?�r�Vf��2	/t�֗���M�놡�YX�4z�X��RT�	HcTrXD�o����p>�t'zIN�wǗ����`�PlZ��@)$�3ٹw� *���O�	�nl����������\m��^����rj}dXD���Ѷ �x{pfs�$�[$i���ݱm��O�Ē��ɔ�����Q�m���'�,��Ճ�����x	ʣ�?JP�y�|wЀ��yڽ5({��q0(��r�ǀ��H�hH�PkC��1�=+���ߋ����[8[ϱ�ttH��#E)�0�G|��= �,W���y����=���}���~Q������*�r�֒$��Zq8�Q�H�\L��e�l���8�"$�5�ހ�������f"�����:�o�1',�I|������n���O�%�_+�3�Q����;G�������
!A��d�>��74"O=<���y���ku�'p%�/{JDQ�_NS��8�7_��h�=1y�@�q�w�Z�� �Y>�g�s9��%`�Y���<mYW��P�/Y����T���ҽT�5��
��~�G	A��8��߅_=�4q���]�ϧor���i0�[LU)x1�{��S33���jf��^�6��مȈ�uG���C�/+#K�z5�Տ��K��v�Q����-���������vՕ�R���GU`��ݗ����>�vc1Ak�)o�'�58�I��ͤt]�c{܇��!��4�.H%r'���G�@2����[��o�����۳��
��Y�Y�$��kbt��R��{q� $SU���m���mւ�rr�o�%%p�o���^Xu��4�����z!��[��-��-:%��2���:��=�+�{�h_���B�3��%m� "66�~�\=3���s$�Cb�O7��l�SA�~�׳[����oI�Q�JF?^�Y�����"�6M�\���L��省���y����j��j�d)! ���O}��j�沆������cuEʉ���"�5��|�[�Tnk i?���k��^��o�ς���[&�vg[q��Hh��#�k���MiR4#C�i�-2�EW���	��@w�<�J�h����\%��s�$L[����[y�BO4���u�ws���3���U���@j=�����S�Q�/�223#���&z�y���XH1/I)(�q�»B���#��������ZL+�C�|�)4`f���')�R'���XG>�ծ'p8X��֎|���_z�M�H��}� ��뇕�=�i�T�Y�8V=%�(��g��ZEt�C����ͤa�:�S�G`a\V���pK1/4/O>��8u�W�;ZW�{Pt6�F��}0~7�¦mgxuF��k����+���I�8�NNq��Oc�����eC����n�z��?{��x �\%��z�
�J��ٔ�	�]�*�����`�i�,�dƧ���ؒ��f�ݮ��b���|�#�"�B�1�0���S|D��:Q+&�p�K��J�v�}����Nʫ���/�6�.��pz�ϝL V���{��cw�fׯm�۲ӼO�W�qk�uqm�C#�휭����P����`��-鬟�������+<��8
�����JJf�-U�0���<Pd �&F�}��mr�����D	�~��f8n9������1�V'�n�W�i��UZ�!6��K<s �d(v󎌈�>��YX���u7�P��^6�@�^�>$�B��b�H \�����CCP�!u��E��,�kk��YV;�|�:(TT�	�:��íYaM���'zt�--����q�zh��SB��'�ij�U�?;�׷�+�
��Dh �xJ�-����	r�4��+I�3*�A5|��!��5aDR�H�����~r K2������9����Y���k���XŐӁF �f9|�č��Rvl�e�0/hB�����ID����a�ũ���	Z���S��Sx�V�-62���2�� '�=�4y؏��H�T��_�3�p.�B����4t�z�V���.3��O�]�����Z�I�Ν�¦�4�w��D�B�w$4��'(��j�"�5=�K7�^��$��9���ǾvW�w��ty��E�(U��JGĬx7;1�B����5K��؁����G�`�g��@.�ly"�yJCc�\�yfFoa���|�nD��/�.�F.GQ�&+~�P�:�X��|���j�Wpp���Ы.2$\{1��(9L/U��3.����W��O�+X#��B�*D��S������x&�ge-��n�<5��ǋ�>Zƴ4��Y��L��0��i3�)P���5D�^B��@Ϣ=�Gf�l,�|�.�VbB"*��^�vͅ]~S��?���2��@�f�оѿ{$�e�߇�BC?��k�|�y��[������^�4����Z�0�W�&-Q~_K�U�K���Gcﯛ��M� ��D�4��qr�7�\�^��O���@(��H��쬼D��}�+�$�srq���h)Ҝ�;S�^�,r*�8ON�Ґ���"���{�ѵ�7߬�A%��-#�������\{k����Ɋa� ��`�3ӌ��8��~ro[Ú���bZݣ�����6�>�FYޝ�>�RT{j����Wȁ��!�'� r?��v%�$r���L��F��*�m�z!Q�����7���������(�)��V#.J+oo��B���ӧ#�Q��W�%�ۺ�?�>�����ke�F\||�_���֐�ŚlAK���Hd�Z!oi,"kPX�k�O�������F�
��n�@b���=���J�SĪ�ȭ�����D8���g��(F
9��[�v0}�&�����mё����G?��*Ddk4��(e���3�Hd�f�w�9<�m�PX� U>�;a��Y��ΐL�@6z�H/A���$��K��B�Y/'��W�b�=��R��mR���M����V��Q�ּ�?����0��;��ڧ���~�7�aig�d\_�OC��W��ŗ����n	��Gc���X�����(5~�D�b~&X$65��FWN;�阱|j������QP��f��vr6�/�{�Y e�2g�}Nh���c��G1������z��m���u��4��«��e��z;7N|~������ U�mF��4���Q読��j�A���3J~��t�u� ����(���o/":��#N���
E�T	dNxP����WRP�GO_���MW���{m��X
p��U�O���tq���ɡ}�7�/X�J1A�#�������s�ef��I7�F�u�&þ�c2�sw��������:5���:���O>�(%���Cc�SdF�������Y�D���1ǺR@}#�����JJ����@���d���[M�^(�Sfo?��ini��O�͝\D@EPh;��]��[�_J�Y���\��'O҆��N��q�a���D������u�ua�K�� #�Ao��| ����l�	x�]�W䙶02����Ä�z�-i�F>%6��"�y>r�3�v���(;t��?k~|#�V�5��H��L��8u\_6pR�^9ZU��	؛�,�J��sQ��� [���>Lѩ�&,6����&ѵ�����u�ۦI��l�P}�	Ѱ�M����*eY�nxߪ4�kV�ٚ	B�	 ez���@%��$:����D7��t�nnH+�܈:u�5?j�ĸb���N� �ؓ�?h&!Ē+�7e���B�ofvU�!)� ���f�'q��v�y����PoZ����E��޷� ������ö`�Rt.�q��a����?��8�����|t��|g�g�f^���3Ms�$H�<����D	Q~�=ܼ�C���
m֍�y�e��4��@�)��=��-),�ظ���b�@�B:�cR��w��G!#+��������4O;IX�u2h�_��%�ܖr����=��OMJ��7�y�ɋ�J���Ò��v��6����4ޞ�FA�<s�*;þ/����>���k�R@��p2����'wN�lLC��])Z�`�F4�?wd�^�90� u����m��>�#{�4E#k����&��֗����ﰰ �_�pU)��77#֦�E3e���ð���ŉ	r4�_�z	Ҵ����pd�M��5o����M@��ܱ��(ƨ��H�_T䢬���~�/�/�Ș�2ܔ]k�9���J��-kW���Û�T��rE��>o��J�q��� ���L�UkAj�xziY��I�q�q��vG#��lm��%hy��s5�d�}ҭ����o l����%&Z��0�E���xfvV��*lA�#��Q��`:�	y�e�h��U>�����V mTP�$w�E��-�rj@�Z�(�O�;�Id���֯8d*�ӱ�[TK�waU�_|C��G�]�����1�0)F�J�;��&�c��]�ȑ}��Mr��J2*��d��c����h��"�,2fc\�P���'��<����#����R���&+\��桻dm��kS)�J�����O�s��@��JV�o��>�D/8�������ml���{s����^�p��eD��9�W�u?u��f�tÛ�<�?p�<��y�81����*7�k���rȠ���x���f�3���]�kH���,�r��XJt	��	����������A�e���ɴ�B���Psv!�N�	�DOg=��g�̏�����䒃T�J�f��������x��g��U]��E(��o0�D<q���GF(�F"���2||�Q�r�O� J�D�g���$%{�j9��0�l�c�\Ůէ	`Aً�O9a�YK�.�*7!�KD#�����&��e�3h�إ��r".̾[��EQaa7�w����	6
��K[�At��e�����i�=?Xɚt��᝚�W���ec��ϣ������A/��HJJ�Tļ�޸��"d��=��߁;PO?�I��P��,js-��I��AX�Է�s�.��KJ����oƿ��wz����	��%i̾�� C_��hr%(�w��/��4�EE��@A��&�:𷸟����P�k_�t�2�I6�&�۲#���9$+{6!#�;W�󕡭�<T�'X�hX����H5	�$�dL�}�8�F�����q�k�|�:��S��j�h�_hQ�gӻ���@��~${t��������\ah+�`�U�������;��5O	1�q����k�?�D~i�V�}_|K���߇e�|i���XevKmaG�܆�vב���<��GG�}}�I�R6&i���ڶ���:�y`����@�A�@g)2��lo��2W��qUm�X�o2�b�h��.ہ�R��>G���
���#�~��}R$K6�am@sc>�*Ж�OM��7��(�I&7T����X]-=2�	KQ���쥆n�GZ�q$v��$4�1ęu��R^��G�c ���sB3�{Cպ�n1	�X��N�}�%��L.�q>��b����N0�����lY��ɨ����e�^G|����c��E�n_(��aUb_�"�R=	����fc�O�f��34�FmHc[]ň���QKMyz:>.9�=���8�>|Q�P�7��U{�-}gb�{��nM[񊹻�K|{<Y���#�����oT�q�MO3�S؂�J��$`�����]19>R�c��`�L}����,�`�'�/�#+��G����^4>mfDf�5�.g���Œ"h]E�l�OE����f�5aqP$,�j �6úc����S�Y:6)������<I�o�;9:����4�!�WC8�f���?/i�ˤwG�Y��Tq�/`0�s�=_)߳����i煱2��oi�s�@���G<e�	|Y����}�r��`��MWW���z	�ck^n*+SSR�|�
T���Ǎ'/4x��^����O�t~�|V�q���ɞ�q+9�*�a����Gl�������!��=�fW����@�c)y9n�N�u/�0@� �G7�|��m������QǺ�k�Ƽ���B)� ���Lѫ��Xc_�g�0��fY��|)�&��w���3;v�p�*�p�^m!�,��J�]o:�����Xw�l/�Ј��� �y�>�N�ƕuk�%�S8MAs��{�Yf�WNBП��������KSb��^���M��MO�Ɂ��ŝ}�?�����H5G���$+:ÿ��P6���Dr�2z��ѐBw0���A(a�\ ��V��c]*���/��:	�b:%��t$�s�x둝����\�;�U��G���߁��y�������!�'7�\��fh#Q[��ve��j�!ܦc�h�ʲG��D��	�����)]I»\��������`��ә��nړY߾ 0�96i����I�R���tE ҥ�� 4T�a[�+XR� �(IѲ��㣵����8����"�e��C-��5���e3l�k�Muj4�����cy97tcek�I4O.3ytOէO�w(	�$$>]y��91IIa������P��tшA�c##jNb�+c	�ˀV]���|��^�S"�� y�`=S�z�w�_�٩��</u�B�)�K�2K=��'n0���:�:��.8��"�΃���f:�j@n���?P�L��H�����C[[�w�<24��'�D��2��xY׮&�xD"ɝ�%�;67~A�̠%�=��y�8���I��Iu764tLֻ�B}��Ы�A3���@�,��pȊ��Y��DƣǏ�
Y��m��댾_��Yɦ��r�^g!��T����265�Ao[���4�iD.�t�O�(P������C�RN��#�~�Z����4�$�P�o�V"���m�"`rg÷bw��1��!�-u:Z͵��#�/#1��{f������I/0���5�qm|u�K&��_�� ���?�E�����A�.�Zk��ң�#�`�)�YC�6����5�>4����x����,66��"�B*�Ĥ��+"��Oq����t����t�%���7� "	a�MEZ���!���T�5)$���=��10��z���Nߥ�����tm�֪����p�Yォ(_����^v�ڄh��ީ�:�EІw���pQ�������*>�|�߶ߍ��FT���5X<���H�`���J�k����?:~ed<��Y�%��?0�3ߤ��rlL�0�yt���������] �?j�|[�w&6I�,Щ�g�O�dH���0�)O�)>��0�����g��8p5DRC������3�:x�h�/p����aqnBC?� �ߊ�/z��~ YJ��J�����:��u�#"���<�.K�(��cZMI�Lc�ZN\[AT嵭����
,C��<=��c�{��xn&9o.7u�2BY���\4�����?_`#�ɑH�cBa�^QwZ��3[r?:_��*�1�<��f�7g�}�k`YRn�����{lB�1�m�.�w�L��l�h��9�V�@���
[�a����lƸ�����G؛��楒�]\2���4�4H���-%��_�񃢑���"riO�bJ}޻9��S`�<�ώӞyy�$����A	�i��=%v�v(�S����]f�ꊡ�2�޳gϢX%���t����*�\\����p5-X���s���^`P�,}T��fZ�)�x��������qz�x�5pS��|��1��������� %C�	: ^�v9������=��l2��--�2����칛�y����C��Q~\}���ǚ�9<����t���������q����h�>������1|��
���^� *x�T���D+�M��^ sO����������(���j��k��{JM��@] �d������ma���XX�;�;������A�]��r ,�oơ�(��T�?��`7�+6������1A'Z	�M�G&��2!��{û�K�^M��u�v7%�+�gk�����]�ul�z=��Mz�R�v�<Ffzu5�w���>̴�N[��D*�c}=����%yk *gs
��\_w�^#�����Au�io7fNN��K2Y$��"���PM��k� נK���N�+�	�-��M>dުC�tDP&��餫�¨=B��ˣD�Ք��'���>��ݓP��P�]�]��Cm��kfC$Wm��c���(�q�z�o"�ڍ�<������l��Au� �aSkJ�Xaaủ�cyc+#ǁ�;[�e��h0Y:���Ι��d�7����"ꊇ��)�[�R<��3��ܙ��\�:����o�r6�A���n�����}�t<��'���
�hܮ��������g+P��x�5/ҚL����,�s��cwH7/�Ytd��0T`oH�b�|^�4O�\�N%�J��<���G{�\Z�6sMU��6n+����N"VPK�l{v���ɶN*�_1^.��(+J&)�kɪ����;�������n�qA9�p��]E�Ũ����⏬��}4�R����wa!!����5��@�h��E��z�A�E�3wnj4���L�Q�b�?��ገP#��D�g���w?v���y+BR������uT���Ń�X%_,��������3�v��?����h�N���Ŷ��1���p7/���NP�B���5�#�WQN��D��ߜ���2�B��y-�����'zT&h{ěۤ�r�N�-k4����y�[� � 1~�/�7ʾPc㪴}��"H��R��A^Us��.G"�^ ��=�:#�	��uV�Þ�2�T~�t��簳,�0�d��uLE�F�F�[���wI�(�(�����r��� �F�u��he:k��8�O25/!KN3�{�n���>2K�g���|ӿS-������1�^��6wת^�M��>�O�^k��,=��i��Ͼ��}?�H�@�~����GxW�����2�hr#{�1�)���^I�<Ylm���fXN!&��"�����Τx�=u�%.�9�k�Q����Qd���C���F�r�����Ų��>Ǌ�[�e2�����D��]s�,I��W~��Hw��7�����)$@�0�)�TF�����[
!�}���F�N	���R����tO���waŶ��"I�:Pu6�w���p���>��l8+��M�*�+=+9�i~-����;��Bf^2�a�%������V���iNS�9�i��ޞ����Z�x�"�IKQ�e��M�͆���1�ԮEnb�yЩU3x����HZ�ظ�,�n�d�FE��E�v�V��IC��T ����l���O}��7���Z�N�x��W��8�k{v!�<_8����wP)�C;��BT�P�Z-���ocǵ�ܓ3NJ�=��7�p��D��V~�,	���w,Z�����{0/�O낱|��������<{6G��	&��(f�������6�C�ze��H�%�FR"< ������A[��b���U��7���j�y�����ꌨ���n�z�!E;~�/)�e�������|��y���,��ȭ��$~k��w���h������zM�H�^�H\yH�gU�UX8J�i�:�lH�do�r����/�F�.��s�_�wͿ��7��:�v�c��i�4�O�#��~�?���](%~:���#t�w��;��]܄�K���#/�4.ѿ��Fq#U�[W8�����5Qq�}��M/'�1t�l����g�wN�#����vv�3�"Vӓ���/+F7㙤�I��x�����K�[9�����,>B������3�3m��f��;����W��:{� OV��k�z�O��Z�j���� 0QK�I�#�+&��όX2����70x��YnҸ�J0Yz���қ�a4�C[�.�;*��'�A"de8(2 �($�nOk h�'���t�P:�����₠/FO�M��s���)��6����eNsN���H�+����t �Un�{���4��[�u�o � <�����Կr�/ٰ"%#��ޏk�`Mo��ӀO�Bwq�,�����"�s�-ػ��赜�MA�J&�d	I`8�X��ӗ�1��5�p6}�0t�`�ÎO�7R�#}�(����K�(Ⱦ��
ߴut$���'�,�FWXD���e{��}�v ��ᆔ�L�@�����B\l\�����֡����q}}}u��hccc�'����˽}}Y<I�s;��p*���8��,�%R�D-�;� ��i>�5��@��Nwx:��J��772�����B�xS[�����$�3��_H�t�&p�y?��Rґ��qo��~m4�y��#}̨@�S��PB�]dn�q6���)��� ���x�iF���<#�C���2�_��W�'���2�����W�t�ᓌ��LNN��>���b��[��YjF��-�V���զ��t��k��i�s�*�6�r���Śbz@oN��
8�T@k&��d�j��XN8GwB.�>-���umb
;
�,�:bSJ}�֡=�;�+��0�Ww�T%�*ec���}�!���Df���[���/�3R��9���W�vu�:����ۋ@�N#Z�fڂ�4<�q֔����|��*�QP`5	���Ҿl&H�ΐѕ�J��Z��'x��]'��(0��Ug)�A�=�n%����D_!+������0-U���N�E��,̥��L{s�?�9����tm89e�Z��5!%�,!�<�dl��b�X������u��^ǳV��w����X��c�'j5X쫙�����?^;C��䣷�W�x�o-����(_JA�f�����a�`Rؘ����ޖa�־�!�X��:�`���R�*�jEB��5�I�6"��n�x���7g�,CB��&��*��X��##���+82��MI����`F�'���nQK�,G�z8q���D��7t�-�v����űc���}�(�7n��R�#���o`�>imj?�����y�d��T�̵�~��y�J��g%z��^��J S�C^�9Z�~$��"��2�1w`te,��Q�Va�3�a�x�3X%��}r2iU#{��&��>$�C�cza�����ǁ��7��
jV��S�X)	�lY���;�K��
ᔕ����s���p~I��X��mk�vP��20@�������P3u�?���.nQ ��I��Hcy&��	:;"2���փX��ӧ�u���r,-��r�\��cS Y9�"����1��J��7�'7��������Ve]۶q*jB�@�|��*ҋ�r#����%h���\2���� 2Z�ɵDi׿@'��Q��¹�lYkW]3�c�����'w�Ѩ5/�Ҿ���G>U��;�J<�^��RcKӗM&��Д�Ԃv��>�/kJ��eΤD{M9�&�~,/!�T����/��`4q�p]��R��o��J���gn:�:D�(�=����C���&Ly�Id�����^��O��$�f�hL��}k��=W�,)\�	lT �db�%Qw�{\�|�=�s"�4����Q=?z3��Dz ��GC�6���K9k�6d���wH�c>��$ߒ>s@�OMA	�^�h䫮&#Ŗ�����~/i5
������W8G���pI5�����<E�i-"ݶ6Ҡ��E�wˮDV�Û�ßX�p?��K�4���]�5��-F~�mF��G#5<�ڂ��b�#)���-s� ��Y���o:���5�J��iSG�b	��D�u�Hd�`�#c�bz��޴*����Y掩)�E�:��A�pF	O����L���==�P�!�����$@R�L���TdUӟ��L�f�H�ݞ�ꩍt�^��(C�p�;�W�`
�Q ��3�C�U@���[��tK��'�n���&j��sGDH�ކ]�v����p��N�$�;�Ǚ�\_7��N��&40�S�R�Ew��-�`�^8�|�~�Att�H�����r���ǖ�-��-5����iz�e7����JY�r0=?{�#	�EU|�=����H��wz�MC�m�a����!��v��3ц'�v�M$�R#�<I��M�	߬>^v+wqt���������/�|��XX�.JS�e���@ݱ ����hAV̻T�P�l��.q:,|TY�����ܕE�N����)R���{�=��5�W%�n?�)QZ�����}��m�'�NQVv����ݦ�蕍XE��\	���<��k;m��4� ��]YbɄ�盽B��l1a���J�R�E����dx�[�i���%B��V�)��G���ל�.�g~�e9�xIH_��}��d�__�"v�Fu�#�X8��q��w\LU�����G��1Ҙd�\��F_@p%Y��x���k(��Qy�8kr��	�)��7S[݉7�]aʟ$2���P�5���Pu��T���?""�ұ�U�8٣8�3#9��(�H������22BV6�J��3�w����?~�[�ԍӹ���|<��u]�Wγ�ַ�<ob'�vF+� �m�<�k���R��@ʝ�:����"\Cګs�7r�X���*C.6�fN�� y��l}�:�IO�S�2o����R��F!��ռ��Q@F⊐�u9#��F���hV�h.�K
0Y����V�)�V5�_����%��O��3t͏t��q<ڪY=��c�#��-��gX1���V��w��P��2�����+Ȼ�z�	�>벢��z�����[��I�3��{@{څF��\�(�I���y����VYuh�����8��l����J�Zg+^��_X�1��_= �
2~�D��b�A|�̢�[�յv�$)�ӬXOㆉx<w��e��)�4+��e������W���uiV���[&u���Ra�=,{(���'jl�Qe���kn� �������%ý�%�t�ЙtޘC�ﰹ�z�,#ic�73�u*��e�-Йtv�!ǝ�q]8I��L�F��v�ߑ��y��C�E�����6�P����4�Y��W����)",��L��t�Y?��[!�$����y�s�8��Wj�]���6�њ���RKU6zѫ.e�)}�M���ڕs��X��/�;}� V������m�߿�KN�=緍Cb/�fЍ�D�_I}x��K��J�i�y���tŘ�dt����)�S�*f�G�-܄���P�^+�u�o ��;��X�$������#W�-�$�����͹�\���;.���ƺV��٬����z�/����"��4*����$լ[n�X��h����Ak��F�?KV�!�q'1���P�+��*C�"��r�6�����2Z�� {�cc��s!V�OB?h�1��I/�#��}d3�/g�`3��N�-��;ԏ�N.��E��a �$k�t���R>���Y��1�2}X�W��z�&A���ѯ������tҴsmOr�fi+V�^�B"r���ik�ZHɩ]*���;#�~�GS`�swY-;mHd���L��d���n5�Z��=[[(벛y�>,,�X%]��q����[y����irE���ٽc���9��hJ¿ou��b�Ƴ�m�c�
��z.V$��~�D���Q�(�F+��y\
H�X3����{0��p�Ha�snW���h7���	G��Ɍ�0hJ!
j{��_}D���f�<��f
�V�s�E�<��u/^�3��o����:u�}�����U��ޑߏ��t-�+�=�'�ҿ������d;-����n�9:�yR�뗗��Dk�+�ѧ�+$#���D$�j�Я)7���dYu��nq����W�A�VF�-+���cP/���9;\�S%j���|���&�Y�?�X�O3a���'ߗ�I�057o����6e����}�n�JnM�� ZG�	T�/�Ɍx�F�3�4�fOڀq�(n���#�5<��$�F�k��~��+iLV�W�����V\;�)K{:;-����z� ���`��QF��u��3 ������ɝ�o�$����t���d�'hTX��nI���δ��� ���]�����GT���O7���M���5�|3����; ��<)�S��{���u�2��nթ�l	�����s��|��&��T��;����j���L����ҫ/�2���	�ͭ&R �����+#��x�e����ڢK0͊�b����T��h�K+PI��S�4�׀|�)���"�m/1�H�`��%�>�_�㭮hg�I��klW��I�ۅ`��@�S�ݢC8��N�o���m���L�?�������{!�Ҁ�z����\\:	�q��f%��ȶr���]CP�.���!�0	��&$\6�k� �7up$J�׉��Y�����'�`.�����gS��%�'��2��?�D��N�Y?���H���?;?������m/��G�)��X�ʱϏn��]�b�|)�}��~��E��v٤����c���+��F%#����i����ۮ�!�I<�h���5N\vְ�>D�P�z_���B8%�eM�;�����r2Q=6�0��}	+8x��QGl�`u���NB�͗�	>&˘��A~ͱ��Ԟ���y�X��e�]i�jo�G�[*��-π�a�������4tZ̪��R�-^�����̩y��G���M�B���ʂ�Z}aa�l�w����e�n����'��J�C���H$�TAg^�]�~��5@w���H������w�sN�/�L��"ږ��iپ��z�7����3��^i���H�2�.��aD�t��#�ҟ"��k�4}�E㕡��7PI�
5f�H�G���!�W�/��Hר`g,�������hX�=*������V�hc)�F��_�grgU-����&k�1�{�	$iؽ��3�0i/W/`���r�C�4���A���&� �0���V��3ir۬|�@����Is\o��T���3�6�$�'��rzl�X��8u|��߰��NE}�
�n���2wK�Jt@�+�3\���쯨��IL��w���N�c�O�G����G��Ľ!W����cͭ����+JFn���X�~�W\0����EQZN�20��j`#E�?h��o-�-��DSL�|�J����F,�	����;V�m!���b��}\��fp���ͺ�)�pd�ud�+�c�g/M�e�
�I�Ubo����M��}ۄ��\X(�(���X��g]��]~	����ͳ��KM�iΣ�o��Etު?g�x6��p���E��W�g+7:�;��><3���S!�t�~�p6#bFjj�M����
�Uе[�m��j�>~�حH��߱w�@�6S9}V�c��҇~P��8��e?�2_P��4�[2�y��aB��ƭ���m�D�7H�lJڹ�>}���6H�kƍ�\�X�t��оTފ��ă��6Nt��J���X��M��7I��$���E�T�+����k�%7������~Z�\\���>`�V�P� g�j}��X� ��Q9˒ ujW�y�;�W��B�*�@���`���_Ǯy��2}�h{bD '̵G{l�:Lsp�2EHo���{6Gk�]�d⓻�29�ႋ�{骏>tdg�F,d����:�wչI�z�ϋ��u
��u���uNQ#�SyB1V��!��c���8�j	Ų͍�[�2˒vrw0A�mq����{�^�ƃ��]��.7P:�`{Ȁ��/�my�|
d��߫Y�,l�-���2����!�V���'�.�L�2~���
==υ������ �L<놖�7�ێ�6�$tx����c*A8���!dݒy�)P��#��pI�RAc$�Ї	�Y������&��e�]����LT���<�C܉�R�9�ߘy���^F�'�G �#�ق\|Bm�9�:�ӟ�S7��Ҿ_`�TX�ǡ�~�gc�pE�s�
\Fi�P#�uA�$@y��W��JF`O|�~,�>�Z�����9����2c\��X�r�t�������; �UV	}���H�+�g����z-�����B��I���^1v��ؽ(�=���j&+v��9+�ܫ�[:���$��<�s>f�����?I�߁��vx��7Dk�.��7��}�uI�rל����`�nʛJŒ*_:� y��͂����`��ۼǇ�{z3���Iz�$�yX�ڀV2�sv�	:��=΄���(�M�Mm��B�R�kAb?q�ċ�����3<4#��5�!M�KI��N���.N�����H�	9A���0H�T1�=aX�����v�魼A�?�5�qwQ噤�II�W�x�P���e2�>����XA!2�yW6�/����s�d޽�BZD��*�i�H�S1�1/p�/�
��+����m��;!�V-���b�p�N��*׳���N������P��C�^���O�5��,�->�A���N�x�F�����] �|�τu��K�i��^X�:�e�Tl��,�z����"o/�y3�r�L���.%<r����r����&KM� ��n��S�M̶�ir.v��qmT[h�>�<	���QLi����i���EFYי�0m��ؒ�nJ�(�Z�*_��1 8�*	�&L�X�i[�W��бe�`�>{r���Mi��R�� �K
�*V3崜�1g1�B�{�5��1Z������Ug//��G? r�M�����yjʚܹ�0U�QT�&S�E|y�='���D���?�c��MZ�)��x���q���c�ǼL�;*�n��mn��${԰7�24�XYJ�?%�r�T��2	3�":,�����땒�E�@?��Γ��Qg'^�;V1��z���ݟx��q�T�ʐj�����|Z/��2� ����������P�"yHl2iJ�و�h�:����|�D�@����E���I0��cP�`��ڀ���]��`�q��ɒ�ڞFC�`΁�U��W����m.�ۡ���/iVv�~=i���S�F�03P�83�*�֩���,(�B񬻒�)��Kߍf
&����+z�Rf��fQ��޸���+��Z8����KV?��g˭�f��^ '��ʍ��u�jMѢUb��X�K"������l��:2Q-�StYBNꚺ���A���
J������bx(�����嵲B���9��馐�]�=�^���W���� ��X�%ɒ�U1���.�/�x��!��N��`���Y��E��|�_�Ы�Y���G ���+'A��ȳ+,�*Q{����a{J�ǚ�ux����a��vv+#
���?*q0x>F�i8Z�N=�\���r��`���E�k�+2����%Lt��W�̈́g]��L����.�?Ҋ�4��s�[����hl����[T �O�����1���w�����a�`�����Z��	��\� y���T�g��G~S��ض������/����6(V��w���.�E}�g#��n2�4� Ӆ\�5T�j���;�J�Uk��;9=�J��O%[����_�#d�6��[<'G�j�L����4��+P���z.�`y��"r�9�ED�j�Ɂ�f��Zӷ���=�����0���_\���M��|]�r��2� n�B-]z�U����������#�%�xr�ܘ��whd�OJW]Fy�}&�j�g���R����0{���Ot���9��2���6j�v�_�y��Eͫ��\0�s,�暦�8㳄<؞�]��^`M�2�{����6y��e�nH�]�������ݵ�w�yi�6w�F�@찕]���/w�����,b]��GG��'
�
�yՌFkv�~@� _��>�*���O�ʝьqެ�����^=��`��Wߚ*�v��w;L�l��.�2OA	�9��͈xl�#cc�I�۱�x��>"�<����9G��Vo��O���a5���ӃĴz"��u�ܕ��mDG�k��Q����30YJ����/�}q�5O�x�U�S�R�u�����.H��ѿP�Ԍ��hu�4쯞e��0�Pף�����L���q��h�M�޾4읏lȝ;u�ե��Ti���K�����۔�+?]��!}v�S�rNIXe}�eS{�_�������nwF���<��͋�������e���P�{i�D�{�e_�P�����c=q��;A��9p����z/A2�\����rz�Pc��mRc�|r�ax�Y�"l��w}��Ŧ�m����s��8���v.%�O�F�.��'���E�d���2�v�������K�rZ .�Z&}h9Mw&�������!颹 R
Z�¤�М��Z��(^ �C�/
�g�N���-���f�]Ÿ�uv�=��ec�������˿����Ț%kP��W/���юsT��n�ۀ���fP�����n��J�H�q�u��G~h$��:r� s�����~����3$�Łb-����A�����̿	���׈*w���M��װs;mZo�%j�Y�ԑ�:V�	��J
D�dO?-Y�����jiC"�3cw�|�6��O�/,CY�-X����?����h�������"Ra�����
��"m�%�^��߼q3Yږ�g_	���-�ue�^�TW��dӔ��������8&Id�bA��_�U·����h̃7��H�����=�2�����ꠡ#�uoh2�O��e��0�q	5N��՛آbڬ���9@�h*��}�(*�����O�g=��I)��&M��p��FZ㕉!,c� �X�q�(<��D�~�������nE�t!��fǭ�y�1��q/�,����]?~��bۘ'̿N�]�.����ej�r˰��|	EG�x�؅,=�M�,���\��){&�K��[�;I|.�4�W�H���I	��MM�q"
�8cv92��A�ߒ�v���|5{�'�o�ԩ��x�$��%%v�����!��g`66>�~ν��´�e�b��6�-)��X�1�)![�o���y�=$Ĩ��?���J�d���u^0�����7��)��9ɺ� 8��:/�
WW��r��p�{�MQ�����h�dL�t>�'�����
<P�}��$�ߤ[$�xՂ�E�M��� ��Y���I�.�-3K���Ei�`�-Dy<��RBvnmw�M��E�&���m�(c�z<�w]Uno������>�.뛢M�J�H�v��,��.K8��h컸8P��P1jRV��+��^Mc�˲'A�f2v'�sN��$Ф�?D!>�&�o)ǯ�脗�s\�a�������ܛ���(�|�~&�~�sl-f�=}~J��'������4�4��"��o�=���*�ƨ3��>)�*�f3�汌g��G"���`_i�t�[)��Ő2`�O	���e�A�������A�������Cƅ��s,*IW�x�,��YX���Z�e�새�s�2����@��VAW�e�b[U�A�%gkiI�>��7��:}���^Ún$�*�Ә��7~Pajj�<wh9�o��ɹ�����Qby<Ww}`��0/ҷC�z�;M����(9)�����W4+nXB�쫦ᳫ���#�+��.���➝&�y�A��'�k*������zپ�v{?�����U����jS��ݽ�/�W��7.�Lr�1�����w�G��e����_-
X$fda/�d6g�ͮ`������oy*��hp�u�v�;��n�L�%ʾL��zy��q	>�:�~O�����9�
g��/���a-o�������nb�2����su��"�`!uַ�'Iy2>6�-{"��P����^�N9<wLjh4�M��s�U�"�_��V:G*au�� �*�D\P<O�0cՌ�x_�dо⧭(U�b�w~[�s
���X%�z �齱��H���H�_ׅñ��M!t�yt�ꎽ4�3Bgw�eJ�I+E��,8�p!{�l{�{:���d����@�Nq�s��GG�����u��~�C�=�m�˲�!���L�ǐ>�;��B�NK��ٗ4]c�-$]��א5��,&���ˈ�O�����ޖ�}A[_����%�WW��1c�|��`��W��&T��[ҽ߻=�����}�J')s�<E������K�-�Ejj嚼�Jc�lw�J�߿�����u����&^����5���g�0w�GS�U�;�x��<\�2��
:�����Cc�����f�����Ph^�?c���=/Ӈ�E�A5dZ	<3we��]��t)�!5��r|�[�� 
�_t���.^Ä�V2����j�^+u����O���~Q��I�V�j�g�7|)�;<,���?jNr�b5�^���$����9���d��BU�o��ҋ��dC*<�z)�{�g��H�i ���֍[��
�H�1��U�]܈���l ��CP�6O�-M�[���]�����!�,�c�����A&]CX�vh��_mD�'�f3?�A!��"��T�nN?��V���N�K���He]ψR	������2����Pͨ�$�i	ı�Boy�Q��~`�pA��s�p&|Ȉ"�gHm�O����B٭
�����`ĘZ0 ��VGR��\��>��"�߳�H���g���{��=Lf��'�J���-�����<�@�����2�Ր��뙇}�n�Ή�=��̓�8՜C"�����
�	[	[�{>���"�w�-2���5l��J��|�Ps�g��@���*�֩ss����Ϙ���U��+8N}�{^U%Q�yq>H���xM�r��&��rB ��l���=��5���(N��72�o�3��ٙ�#R~�)w��
���������ζaQ���k�s�E�"��D��`�_��"��(�M����U.,���'� ̀b�������{y�6��i�'���aMz��d$}�FRWv��(U�s��2�	�2=�� O;k~N��.v/HG�Ũ�hN��5S�
�Y@t�AV7� ���lU�;�!�k������<-��E)�� �iƘ���y6�͟o�H���	�nQx�&�wҒ���Rɿ�ɇ]~Z�a%�Fd�k�
sO��<�������=.�kl�;yK=۠��L��}9'��X*�8�T[�:���Ǩv�'^5ə�:�P��D�ǈ�o˖����ʸ����zJz���kͩ�˴�}ח�n����`�>_KIpZ[��9#"��J�F��ee�txϬ���*}#B/�[��L�SjI������L��������-��;���f&$
<�L<����������@X��BR�Ա{��64+��w~B�c���ԓnla�]���1�-�`g�Q�D�)tsJ6R�x3�%f9<�&��6�'�V4���� P�J��>��'r_��)�K�^�w�V����Cܠ��*#�ޔ������A�٧���Ʋ�1�y.����<�3>��Ԉ@U�Ǫ^e�wcZt!�^)���̆s3�����(�|WT�L�~0��$�'�P��13',kTy3��͡UKqe��՜��X����}ʱMp�qsCe�R���s���7���.}6�$s����y�t���(�Ɛ��P*��N�����gF+��Mޛ��ۑ�d#�%����h���2%�4����I�2�>d	����7"�	trk$���ኧy�"�����*9�3��u��H`�6R�MG�c^���܁pE��+W��P1VV[�E�a���}�
��Am�&_Y$�5�2��iE[Nj� *D�/}Cބ�7Jc,N���<�����M2����>�R�Vm�C���]��~�0{\C��x�����s��bR��L�}�G]~�
Oe���jjH{y��x�^� U������N�}�<
n���p�����
e��{qG��\ǩ��3f��#D��"����72C@m��Q]� =^:>�)�L�d��"z9��@|I�b��Ǡ�rH�e�"w��!�l;ZT��[c�ڷ�<Gv�4m�@����DY���i�ЬtG��]���΀��џ#k�,��Bl�r�J@�eWg��G���I�Xq�-^����w��&�����w�P��e� �w�	/+�z߇}Z��J驫�-p���g��U<}�Ue�_s�='(4%F���=�4�����ӄ�3��s�,�3��n����7�B`�D$�n�%�\���L�(�1wV
�_@�~]�#2P7?���O�-�6|��ֿ������p�[�uUU�?]]9	@Y?[9a45guv�"X�/C-'<wT�B�Aa={j�IOs����Pןb EF��j.X����}�I�X�5.���\�GQ����R��v�x��8���Z`4-cQc�ճll��ڨu��x �
9W41'[<����f���U@I�`S�IQ&���Ԓ��&��=���]��|d"�T�Xm��W��Q^�p~�����E/�^�=����9;�����y���2�Z��;���)p0��Q�nK�g���yga�7�6~�ԫN�}-999pj��#r�����q�d��G����#�۷�}�� ��p���O��jLN-3�,b����9j��jz+�v��1oe&M�`�o�e�'��*�N�]O���[��p��%ٙ��3��^���	�R�zn����BH='��~�@���~��ĩ��'�����t��e���^��D�K=d�S��>���,�5�aH�M����NE��`_4�e��L�P�4�Ȗ��k��&G_��Nņ�oH��\�=�&�I���Eڄ}�ѷፃ����8d"�C����{��e�V�Rt��ON�xi{�D*��P7�
1���9�� 3���K�P��ܝ穰 �
Y-?���3x�Ѻ�����7�IT@=�O��;�;�A*�KxÙ�}\�js���9�r�[���L�3���G����2}��E��������?Ɣ���k|��%�-�O�ZU�bp�8���k�I�yq�� =�-�����k����t�rX���-�yJ�2��l�C!H� ʕ���6�Tt
[���=�S9�S��i��>���T����o�e,߇�ډfkqe�BD���3��@)K8T(=\�a�>���a���c=��u�̞�{�_��`���H�2��o�ϵ��dr!_h(�7\%����_��r6�EMW��F�'��9�';�Y_Њ��ٶ:f4�t�֠T_#���t+�f�{�������/5&����,B������j�Ơ2of��d�Bj�,�fn�7�n��1�\��{k�~B�NNŮ�([R�4�s�Kgo5,ԯ�}��-Ɓ��#4�/�7��E)�fvvz���
�T�A��;Uа�]�_���W��\��^Byyy�ؑ��Y��S$��q�������zF�����+ԕ��rP�X�j�k���`~��<�I��_��\��iK,e�����0LXa�]�[$�D��\��h����}ؾ�Ƹ0�)!w?��6�%u~���F��?����W,�����j1�\^�q<�vp�aJ�iAaN��ѪYUR����`�ʻ���5]��!�s4	6o��g�"P��AB�tN h��h�4�FQ���0�|0�3�p��ƣ�0{�~_������U�i��R}(�ޏ1�n9��&q�ı�����K]X�sR�C^��!1�WLb���A	����F��S�Y{0Qi{��Jg	:Z�U��oy��ԉ�ޑ(b�"�%��������>��k�4���l��#c�d��r�V���.���y+����]}�_h�n�KE'�A=H}���<l���%�S�y�ա�&�K�"�J7�kn��y�ȥPŌ�t���o��_6��h���Y S�3��@��`�0�U���Q,�E ���O���x��g�Sl��l""%ޯZ���4������CP��L_w���BZ�.�Z����<ꡟ��[#!�W3�Ս�u X�dx�����a�{��H3��N�PIm��,:�N�X� /�o�_�ξ��hw�Q_"X�-odz�ש���0 �ga�a��<�t�,�\J��Zo��񵪈��-�eNk�$����ZbB��f��K�����d��1�w��C�u��_@Ҩ�	���)T�lEc�d$g��%c���<�m	Wx��.�����O5���U7�|xb'��<��y���0ʤ��#E�z	��װ4���rS'��s�4�Wݧ"�\��D&z��#�V���E�$߇�%��ME}�A���x�� �Ș�vXa��7��p�?*�� �z��X7���e��r�8�[��Ed�Pqb	����I'y��+*�K�N}N�5HOn2�<��|��}��0����C�$&Y����,l(Q��y*f�Ն�P��̟v���WҖO�� R�}���.:�l�%�ܶP��������]4z�|UIEu��?����ΝHYh�C��P��O\&�;V')xv��%�f{��m���M�t�H���,Ȭ�J�%�o'X���#��ny<�%\f�ƌ��q` �[;ڐ^��b�7
������YV`�]�@1pl���޸��m�Zj�e�P���>u��ct��JR�ƣ30��>H��-�2w����h�k7Ϩ�r_,�}��@9��[Af4
�7�D��������7������E�t%EO�T��Ͻ[�a�8��dOGݥB��<��?�f�/�&$͒ݷB!f�����+~Z���*S���?yE�3����W-
ص(�1��Pz�����_ !x�����{[��p�]T������iV�-m#��]j�Ӌg7��T�y.�g���'��!y��E|��N���� ��jE���k��ę`Q����q�,��M��v3���w�_�]��C����}z�{��]�d(w�܃�݃����V�~�ﰈ��u^й�u��0$r�}���o���[:%�`u�~�������Y4�S�
b�m�����8kp����x�����^l�6��^{
\��=j�¯��L��/���rw�>fP��㒺����"xb����գS�آT�KV���=U�ˮ��U�5�3��T����(Ӓ^�t�ъ�(�ɲ���%�4�_?�mZ0�$������$�O5���U�]E�����eM�6����Y*x=T�b�ra\u�v���.K�������*`%M3URP�~��b��������&rW�V�����e8a��T�斷D+�I�/�2x��un���$��v�ZF�^��r]����2WTǲ�@����7��zq}���H�01�,�~EIII�r�j��&���ƲI���yF�Pi�~Ը�,�cy��GK.�fQ�[�n9���B��+�J��C�/�|P�خ�O �+3�ތ'��8��)C�,�� %���϶�54:��1!`��m7%�fZ��i^	}������oV�]A�9J�l�EbF���jp��$I�����G] 39���suc̿`�B_ƻ|�rKO�������0 �N��C�4b�k��3;;;;��q����՘��+�^y䵐>ʩ��XU)ݮ��_�� '�7���D�\���1 ��#�V~`)��iLJ0���m4�X3!�8K
��G�xF139���"�h� a�V��:�ڕ�m�*s�֚?�V��ݾ�?>2�@���I|�:*5|m�mT�����.Z<��k羄�<>���I��\�N&��au��(#ߊ�S��d��n�ܕ-������
��7��u�w���`<���F[i�|e�U�{��H���;|����N�x�=�&{��2�
�L����DUs�~�Pz(���=�K�_u�����o�t��I����CUF����J3�I�N@c���\]�y*ɦ*\��}d_�^��{ �-k��SkwG��C�^ޒVt�Ut�ؤ�6�*�sm���]hèW�Y�ӏZ�����`h�)�����׆g���Ӕ�4N�au�ȕ������p��ka�"ǔ��q��㖐mb��<i�78��:�E_F�Ph�Db~[?�;�N�U����ӧ#P�	�߿�џtL"*]�	�V٩�o"
�[;�m@�������"�� 5鼓���h��<l�Rt��<�}��UWP)@�7�m%x��ѕ���R0V������7¦�j!3�J��M�����G��=��@o�#�@�](�M'ݐ��tB|�Rp�Pts��q�{���r�r�xi�����@M���n�q;�۱z�}j6�����N�����o^������Z�3�M��˓[�Pް�X���*�2�q�y���511�L':�z���N�z�)�ژ��A�Lh̯�X����!חMK�!h�f2��'o�Ki���U78�wZ��!�9���x�
���I�R�O��S&#��a���5�Վ��n��^�Z���&��"�i���*��8�E�_qqqPs���`=��7V����/�� ���B��Ï���{�bf����6V!!eP��Y����jz#��Hy��p��V4���1�Sb���8Qʅon{D�ϯ�a�K��G�Uz���g���Ѐ_�i��J/w-��f2�6OT�:��Mh$����^/�5աzOQ��/t��9������Vw�q���S�D��2�7�P�����O���S*X�	�K��$罬U�h�F��u���L�a(E0o�ʦ�h��ŏ�ϼ_,���U6������Q�� ��Dn\�K�nha��]�H|M���2�tY{����!h����kY:�ae�q�'�B�����:]3�^�.���i�W@}5>��#��������[�E���㽾Y�v��9�~TQu��ZP@�|��Ʃ>�U��
o%����500�8�ĉ���[��V^-�)�*j9�X�)b99J{r�W 4��M����A���
���,G��xF#K�\?�l�^�'��EX����ʄwB}A�@�y1-=���D�,�Ím���w�Ըuf��^ ��0��ݟ���!l�6��Ч��H�x��n���,�L���_O�s-S�[(��At	�ƫ���X�&{j5l��J��t�TI���>=��j7�v`*���l�[0f�G.�%9�l-J��K�����>M�&��AM������?%EQ�`R��� f��4@��c��N��+�'퓯V�akEkK�J�����F��"v~�)� 
���n��㾻!��n-���5r/7��z ���6o�a���8��q�|�ҏ��`��P|o�y�7N��mJ�?{UÖ��^��e��|��#P����
k��#X���˕k��M� v5��S��(0�I�M�z��%i���S��D2�W������-�����Y���N��ʂ�(ɚhM���S���U��N�:rE��r�O�����ȾIy-Ol�LJ����s�Oc�\7�^s�_P��A�W5&OM��r�ܠ�T�z9���g�w��hV~�Ȧ
�9���r��)"�oX\�r
O$s�Ûۘ�NfF�%*QWG)JQm&�t�CoI���!Z)�f���6K}��Է�G&ZL�w}�8㓒 JI�ɓ@��n���/(�O�r1R�s5�76�|��n��x��]d�����G��A�k�P�S�������
c�� N��H�A�{�34��_Zoj%����N[�Ua4+5CD7O�d+��9
�� BO�r�����l����g��?�P��s��o�	g��y���j�M=}m�^)fLk�F��r�!�r4]2��u�[��և�y���j�L�}�����v�EL���l7� �
��ff�>��59�c]�P�Ivc�
b�l��/�Uf�x_J�T���l��J_���9��v�>v�gJ�v�L������$Ұ����"=��r�v�$l�����g"}X�؝��g����1�������K@�Խ�$��eM�gM���Z �&���I���B+��L\m3TC���y�z;8�P#��_�-��Th�Kզ��^
�GQ3A~,����:��9�jA��ż����}[��,a��e������O��M	�9!p���|7V�r����J.����r�����U��S�r��Y����x:�t�sfQ�b��#��h2�������H��54��o��*��4d�= }�u��
[��{NZ�_��(ȘZ����m�<[���׶џ�
�-.ag��;�Q�1��G�d-�1F��(�_�l��X�Qv�%���;h�����Fd��4+*0��B^*��mՏ�T���3T�ZP��R<uN�K ��,)}�iR�0�i����J��[�y���5�����;�/���	��_����ݝ��(<<}�}���F�+G�;�c����� u���|������y+��X���r9��Nh�j�g`8�MnCrpxd�D8��j ��=�XI���3�����^ܗ�ĕT�g�tm �pj\w�YL��!hȦ��[�{Iy����*��(g�|	.!?�z8��;��؉c��$��?�������A�//�I�v���rs����.O�$�l����4cw��2��8qjL?�2��L�ݹ�ǍLl����|�'��$���e"<[�Q��Z|-/+-�%�1�(��m�$�kY�k����OEh�ym��0�B���R����N=�뉶�.��uƅi���p�9'�?��}oM��>q�fR������~|�EG8�r�ߦ�cY��t����Ih�}&��jP]��2��^_.��j>��K��6�+8~���q�(��uEf�a`)5r�<��QW�Cڒ �cTqq�� �FS��/vޓ�m��p�z� ����P#Ҫ[7"��w?�Xx��u�JA���h�t�)#6�
H���3�K��u�R����a�m�����D�U��ՙ�p �7>8��\��tK{J/a��4���_E�dP��=4rZ�Zt�1}����q��>� �!��!O�?#�o��O�V���0�G��e��l�yÂ��f�^�m���RFފ��ips)usD:h�+��T?�L��T\ou��ON���l��h�� }x�P݊��a|[���Fܬ�ɼ���J��y�����y&Dʖ}�2aS(釀-��M)�����xJ���ֹM�H���?Gh�7�c��O��"-�G��e�����=<�t!�p|LT|]A��۽�C�j�o��,�A��D��ā�-���@��>�э�'�V�(��=��#���R��W��m�K�x�j���~��l_�
�N깺s�睠]�`��l��>͢KG�+�_��m����.Ĩ�����{����)=mj�a��OB&����`&�;f֝��� o�NQ3B�c�|���[ ���	�����pO8�x���=;�$u������N� k����4�m�n/G�,��e��Up��Y�T��S�[_L�~���Sj���6�$�z�P����Dl0ەw����V�� ���h��Q"A��LPj?�4��?�4�F���3��c<�#�ſȀf� Vە%�"(~���2���nd[^f�P_�&�u)�jxA�],)W%�đ�d~���nM���NN��WM�=}���0�Dr
#oiݻ��C�Wj�\)��?�������6I�&�k��d��D���Ԅ����j6c��}�����o���!j��/�.1:�{�'X��1�<��3jC���ݔ��uErN=��r�[�ˡ�����Ę�5*Q�k@������O���*GBd3y��˲�>�΄��q��cPe*�]���0�-Ķ�P��[^���t��{f����^���m߭�KJ�d�.�+e���h]p0�5�({꣈V�ʓx�r�X�"Ů���K����hn�ո�vi+�vL�X�.K����'�d)��:�ޫ0�������?9dS��ɮ�tdD�讄�d���SVG����EQ�l99Ƒ��BV��d�C���]o���{<�'�^�k<���N��2�g~ӯh�qiNx��R�g$��>��$��37�#XMuIa�M}�Y�^mB���Yy�~K�ːӔ��?� x��,Z���{�XjA3u��ro���{���F�T��(�<�m��}���i+?���:����n���k�v���B�����0���o�,��B��`�=-�;v��ș�e��m^���-�Њ߶�z���jAȟ1���c�OoN��� �i�q3_e�0q��L���ֲ:��%���������},@�z���%|�gpp�kx8k�+A�4Aڠ1Y'Nݼ�����=%<'*T(44t�m��Z�s�q&��	v�ƺ��p7JN��9 k�Ue%{(��� �t�Q=R�6������q�F���� ەo�ׯ��jjj�_}&�8��օ͗A���33-w9��'vT�~5U�q+mK�':��G;h��J��=��m��)^++ny^��M�����KZO0��s-n�ЃNyq�"K���_g��F
VPWW��q� ��03Lޓ��u�EԚ�u.W�Z
j��OS�Z�0�jLLX=nk}=8��u����2��������wɑ'^�|��e����=�%txE'�<�%�5���S5�����Ur���nCӱ�A~▽VXQ5q�0��sm'"x��˃�z�+����H��X�nl<���}a�޳ۥ��y��l|Rj��Kv���k�ќ�S��a~N��-}��:\37�X�#�)?=n�ٮ��p�F��+}�J��7&�i�􅋕Y�Ž�ѐzd�z%� 6��U��Ǧ��iȧ?�7���I���Sտ�C�9jUA˼{��j�%�Ec`_?u����@�7��"�h�!����'� ��$rL����#ZI�^����JW�N�a��4>8��W��A��'i���NL0ϖ����b�j97�e�b�L�����|о���(]"��S���p~��ku�]%%Ogg��С��̱�Dm��Pm7���{��W<�OM1��Jc^��$���ʲ�'��g����s�R�!����!�&�G��j^I��O���b*��ia��ӳ�f�%v_Yʟ��Y�Y�q��u��ͼ�b��]O�ۭ.s�6�555��v�h��\/��EEY
�m�`}G��'Y����72��yE��8m����=&��x� o.pM����P��ɦ��Bp:o���(]����w?@II��zr�I��tD���/)��+�}���}*�49Z���]���(��w������lV�`�A#%ޯx�����UE��N����Ӑv�=c��J���H��+�����D�Qć�⯛����C�I���J�x�z���>�V=X�#cxK��XS�
��3��RN��`���NE�U>�F�9�l�)֎%���Byu��*PVl��ȕϚ�z�h�c������'%����	�F�`?3���e�p�c���5�ϲ�z�x��2Tߨ(�>��������+?���k��S�E?Qǈ�V81���!9��z��v����z����ыd�2)j넄��L�g��h��
5��i"�o*d]b�N�!G�Dd_��x�	Ý�;����$m׭�	{�VZ^~�2F�� �|`&�yM�N�Q.4�^%_�F�7x�x\��/}��_Y��W��b.�[n��R���]��(��瘖�h�~/�w��g�=Ŏ����?��������,��OM��H���f�)���m�Ճ�|���Cᒔ�]�����6=+.Zb�G:�F��_#��. �C����x�f��9i��9]H1	��?�������1��=�> �PȞ�*IЗ	\H��{�cm+I���	)��'骺��UUn>�~qXwyk������������Fp�]�	i�r�Y��-�Я��x͟�������t�dW��qT�� �ɷ[�J+** ��~TĒ��K��7��D��Ԡ`kk�ãzb���`SsklD�[�34n��l���O���O=��l>��q����g+mi�d�jƏ
�>��u#�~���'�˴���@�ͪRc�=Z���������_�ml��,wz�E�`'C�&o�A��p3�f!�h����?`4^����'���iR�Q$ԭ����&v�+^ԫI�颉�Q�0r����>炶�	y����a��΃lD�)� �2�&�o1��2Ÿc�ֿښ}��(Q ,3��ۛi-�# G���)����Q�V���M��Y��Rl��v�==�Ū�K�A{=���0�*-t:���,U\.�H���a߉�J���"&/�Y�u8ꘙ`2%�?;��F۵�X(�,��t���QV\L�� ��W3h;��í��W��`�w�$�u����@Z^~S��9Y6��Ca������+L���f_�L�W�c{V���ܳ��&��

�֏����&�ߓ�X�������'�/����T�ѻ�G��f[��.'�/6 a����M���i��Vud�}a�;��&ݣ��зdt��|3��	�am,�%�P�=4����vS�o���ʰ��j���85a�@_��֦�&��m�ǩ����X��[iVb^�Q��
���hN@r\i��d�5�_�S������C3�����i}]+56�B��z/�k�]фl����OV�:��\5a���ړ��l��0��0�B�0�_JyM�@�qz%=�JF����vpx1��E��s�F�qvmD&P(7$��R�	h==K��~S�Ԫ�m�f� ���J�9,�����_���S���vW�R��׫5�$e�t���񲲱au2���?X���$�<_����h7^O96�42RN�iS� �D��3D�K#n�f��0�[����ֱ����wA����y��>�'����#0��$�������r<q*�>�2�GX�M�/n�>0O=-gQ�}�ڵk���Wն	@�$��Ss��2^��f�[bp�*5�F6vr.���e��<�u�H֒	���f����e��Q����TK�09�<7�^x���ԯ�ȫ���	�_����6~�Hz+���A`;6":�7��8��e�����YZ���[֨y�r�~��o/a��U(�O�y��7�ۏr#oHE��Q��6喅97A���k�N�@<��i���8b�_�����F���>" S�K�G����/��<�8s�!$�Ԉ��#2�~���;��ȾT(��i���+�#�0�T�2;q+`�����ܜh��r|��4�?؀%b��$tv�$&�͘���uԛ���ܸ}�v��[b��|&,
���Q�|��sk�7����2�?�йq����ʕ��6"a8fO���E��.���F(6���j(;�f�$n���aᎵ]yU�b�L}�-��,�Аkn����"��+�.��*��u���3�U��?�ؚ�32p�[��r���b>��R&�<Y�P��G��[�O#r��J7�^�3�pJ�/Mоw��%EE�����͟{~�2͟���6X�+��)��nl�Xm��E����j��K�h�dLFj%j�4��������13ށ�`��`����"%����҇;&�Px�_��V�?x-����W�� =rn����NQ�A�}	���aGBr97ʁئ�A_Y��iKȐTza����Ċ{�l k�*nO)�����a8nLHz��-�]^�vw�F�tPj�r��۰I> Zzꑍ����!lp�V9��*�؍� ) ��z頋�N=>�U�8]t�od�sq`�ݲ��7u�����;_k^	l�,��˃�tuoFV; q@��p7Z�����l>��>���0^�U1 }v�W[�s"Ƿo����w�`�����f���l��ӣ��1��	nA;V�nx�R5x7�������ܬ2ʽ �5�Ǽj��dۻ�a+�U/�C���Wf�Kʦ��I��N�e�=Ы�֏�.��>'}�Nl�A q����θ��&�B�w_�	W�"ޡ,&���|� �bs���gI�߸0P��R���&V&�c__@Ӡ�+9p���0��+�?N��S�������2C�ih�ӑ#l�7�n����c@������� 2��v1��Er�S"��%�
h"3��5��y纴��L(�O�ssHC�w���2�?�;dWZ��ðy�d`���%4D/��#�3(�)�%��M(]@U��]/����X�xAB[�kVV?�5�Q���b����
�
ac���4��I��Nzaha暎A��IX˱��}b�6�z��qn�0��<7��4.��H��0�}D=��R��7�
�^ �U,�=�m�m���������K���OT�Q[�k{�5�qP^Y���-u�[.�F������[in��Y6q�zdfhtD�����SH�_g�7�,�gJI�/^�|5&�`�����Lk{���_�0�2i��eI�vl���tU�GIc~�`O�Y�����p6@E�C�����C�S�]p����(`v�H���jLM���N�iY":��s���3a��i��_=�*�7\\��Ҷ���,��#������I�9Ɩw��l�VSgN���?�z�87D9�#]#�g3�e�+��B5���^l����n�_��X��f&���ي�o"N�e��0�����8$��}��y�Y�d��=,��e���vb̍�0�S^K`eR�\�~o���F��9�g�B�#�pz��<񔀂"P���~j19-�P74�n$�^�\�s�����--iZV�AbY-�4~3b7.z(s���ׁ:���+�R3`'X�ĚFG_������/;��4��ɖV��Y�6��ne�V%8��C���[W��ސ�X��T�&gg�� M��TVT|ו#P�"�N�ƕs>�%��Y L+)YH-���T�i��X�\��ȥqeA.b��n��E&nE�1�K�[�Xoؤy�X��jKQx1��NSS+(��ƹ��v��S}��n����RPRB/��J���t^��x�����Ye��Ҕ=}�^��ުl�(��NVfwK���@�z$.T(Џ�a���>(���uh1'�2_tm��P?������/<3��}�Fh@}ϕ�������Ձ=��:;��OҊ���I�
3g�1UW����8K�89����]���L\����|Lo}8(&�}c Ia��*.����n��u�R����vjMxhh:�QA�u�����{�P!&��5�vևրQ=|������xs �� 5��k�}O����Tu����S����ӫ��t	� w�t�t�[5��{3�ޚjSc�P��E�2��΍)��f�Wi�!�ӏS�l�cx����_�ul��O����?[ݍڞ�db���T�G�G���Ɪ��w��vWߍ��H�s{e�s�$drf�z`��u^I���j�;��bb���������7��45e�Z;#(���K�f�����{�c��#�/��ޮ�P���%��ƲR���V�(�����y3֜��s��H�Ϯ�n�d�92�_�~��s�'Q��G�[g��ԋio��{j����˳��:1�̙�-��d�v)���f�-�WJ
����:iђ`����tǽ�ິ�Sd��U�����2H��M���1P��Ir�SiZ���r��r���ai��#�j{%���Q�t���Co�H<}Z��6<��vW���,*�>x��2!�������C�+���;�m�˹���6�B�߮q�m�j^+'�g[����/�z��@N,M3�QO�Ac��>/"4�p\��p���"���~0�c�W��cg~�LVĆn��\�^��Z��9���ڍ�g�Oas|
����Yp<�A�9>Å�&�{�c�gN��h�~p3�����+=�a���̓;����a4����z�7Htwt!{����{�]n��F������kc��Z��c^ ��\ �1lm��C��\�	��k�=��`i��~*�T��5�Lpx�F��V��5J�p��\��\8��=8�}DP��(XN"}�:��6������Lq�e���r)Z�z�}�=u!΁���J�|~��ծ�����F_d���w�P�2kl@�v�YE�N�E�Lp:�ʸ��6�x�?5׻]���U�+�~[��&�X|�i��JoyL�p����{�O\�(��XD����1���?��uߘ���.���%���KHye��}]��xYi�(����NǶ�R/�nd�|@3� 3�z�M����J�Z��9���H�0- )��S��4���O+9P<Ի��À:gA�O>v�����������L6+~j������'w!�c��W��C�7������\�N��0ڍl"�#O�f�CY����a���d����~T�q�vy^]�m*����Nݵ�"�jS�T�LM�lO�SeUϬ�/>M��ٺ�.��׵�m�������u�YW`���!��f�BBDGL��0�^���)'���k
��<!ٞ����D|E���u�&�|�%f)h#���[=��,���!%�e�`�{�Km��0��u�3g1�25f�1>���h�ދɛ��y�Wd���%ج;6�q/�:y�	�N������֝�(�c��{Fx]��x��N�lI�<���,�YZX!��n޻����U���cS��M������{*P����N	����v���(�a�W?t��9�Q��,���W�������9�GZ�m�KD�M���!�t�lRg�݆��<%Eˊ禧
��wK��/T�v��i���z�*�n/u�,�����;�Ζ���>�hi2B�_
�J�[���Қ���?\)�s�,�u��![>t�ݘ�.�1P�E7��Q���A4�לk��7B���<H�%w���A�-Iy��H L.��:�\�M,�l��)b�;nm�jH�wePÎb �Z�Y��@����ҳkՍ��������:o�]�M��e.��Y��	�B��5
7���'�m$9?��~]^&<?ϢQQ�J����Klu��8ۭ�xD�.A?�c�{�@��WF$7���m��Ŀ=��g�������rU0fĔ׵��*����8r����yv�gU���u�'����V	�a��\.�do�����<�V�|!$&�U&\��qA�W�^���忱x���!�����΋��a_U������v�'�\<1sJ}8|-'��Q��ߐ�2�))lA����v�_'E#kj�SQ�/�Gb?�x�4s�w�
R�eqrph�%��s�j��g�_Oˡ��+����7�x���Q����#���URY����C����{��ث1�X�-! :�n���SU�V����u^�Q�,LCj��M6�G[B�j������ݏ��h�x4������n��R.]�q4f��׍��3�,���fM7%rX�J��s%&�;��]��H��+)a�]�a�Ar��ʏd�zZ�f0;LEM���=�c����� +�Ia[��d�O�����<�4�&r�ˆ��x��Z{���$W��
��Vv��B��ͻ/9c�ٻ�����#�'i�8ɫ~�����JOǙj��E�'�����řN��N�`�>��ؑJ�b:�[��;0�Uֆ�84S!T��u�XVTR����k},*p+��S��s����n��Q[q��\+'Rj��@���>����g,�J�%�
�Ŝ35�t=M���,�e"M@Z��;�+hik$�l����l|։{|�}��`�o�joK�Ӯ>�wX9K����QN�$B���ѓ�a������[A?��b���2)���:�C^�%��	ti��W)�m4�J111^��GX￧J�Ȳv��>�T��AWW� 6J655a���|������z�nd�M?�R\�	�����?t�N��Y,..�y�pa�
�����5'�����3��� >o�)uzĞ����E��~���;�βݗ��Č܋�q��LfG*�>�	�����w������&-��%�,��P�?p����ń�W��K몧"Y��g{y��Ps8쐙KLa�7CCM�@ch�+�o��-lSB�u��F��m���w��YEf��K����I��?��\��k��_���۞&���/��������;n]��D��Ǽ��3��ǂ%�<��&@W@�U۱v�kR� 뎮�������#�H�� ��aq�Px��X,��' ��͏fCa���G��B�3��~�e��&�����.�w�p�W�a�XE��}'B��'�p΅��F�W<�ǣ��u�	��Ӵ,E�T�IK�|隋��չo6����GHK�r4�P_Nq��RMC��~`���}�����sU���fl�:��7���ފ#�+��N�
tH���C��|�B�GOlWW�ng�
> ����Ü���>�j��#�HDw)��k�FK���1�|å_1����iPc$%r��Ng��+�r�<��F">Kv&�E�$BS���jv<���N�	`A��-�kE�Va��b�[2�u��Qx��/�ѩmv����I?]���ƤB�,b/�\�bJ<r^Q�(������.��Gi����4������t�0�2]ӵ[�����6��n��������s��?3��!-�i�G�Q�3�D�۬|�7����0���Mi�[�Iy<�,�S$�O�F���	�9���LWV�d�-��[ ��GOZ`��w�4)�y�\7EHk%m�2;�=�ug}RZs䯳}+�程�
��C�7H�jl�J����X�'�Ѻ4'�LN�(�ܯC��/,77~��E#5D�~2����.�b��!�t�f��F	TUlJ�*��Sb�ώ���f�m�i�A�КNX�U�9���'�Ze�}�/e�BM�u�[�d�dj.wG�MԾ2��>/V�J8�K�������CZ�^[��*\$�#���3�ϩ\j��_)N���ש������WYe�8����k��Z�����NZ��V�������	I��6��v�L�]�C�v���S#��7���8�`x{[�;n� ��>�� 73c⦟�g'��Θ����X���S uY:\�&���iݫ����J���!��[���S����џ�_�u�����Ɗ��`Z���D8��	���1�[���ڽ�ne��0ioY(����.+�t��Sct��[���}ԅ�V��qa�X��{Vw��oUX�8�bX|�r�e.����y���n?M8|������V[��=�d,�ޯ+@��?1�,�s4M�A/��9s�4#���WEA!ܾU�A�r|����:����/�	{dʽ	�8���:��)�*�*��g�SS$�{@�c2=h���h�|���VR�B�0?���ز���wa����7>��<�.�6';"����a�\�m�n���OL:b6�0���lJ���5�����ޞqįD��6K�/l&D��)����:��0��~G�4���|t��m�w�g�.�B�;h�  96M�S4���cy�1��L���a��GG��CI8t�����FM�r:@9����wV�p����'�لL3�B��lӂ�5��I�Y^|���� �Č)�f�u�ߟ�̬�;���%+���)����9}�wy����0�`�9�9��F:�K5��zIfKb<Xq��H�٘���Y���q$�m�+�e�?9�Z̟�9�PB;k&��r<�CĆ��Ѝ��[�&�2��.�Z���;��`;�sO���7]~ͬ=�[X9Zמ9޺�(���)(`b�ګ�~�KryUPקE��!���1��I	��I����d�#�v�H�ॴ���"\��q�� *~=xS�:tb>�ku7�M���D�u��?c��[������>��A�1mZ�X~�-��5�Wt��8Q0�����ҷ��'�����?�H$)5_k�on(3��:�Ǩ�!��b�jo�-�3��u|~vl���mf��X�6���o�f��d��S�Ҟ9������l�Gi��oi� ����an�+j@Q���iH��zV]~�EN��B�Oݺ����cz�H�@��I�O,,K+x�{��"��ne	�����6�*8�+^ـ�S+9��$�ZgA�3�����J�.VR�v��9�.�R_R���R�A�uj��D��>F�TW7?���q%��o8e�1��}�G}e%:� <B���y�L`n������~�Q$�Uۇ�w�P@�Ը:ܩ�����(����J����aFc�!9Po[S�p���Bܖ�4ŕ{�1!/�+L�����Ջ�:q���V�T��&��&��g��U���ׄ����������g�u#S��*�@7)[�݀�~f�ObE��(��h��y;}4П��+��o�3s)6GA��������̄)�6�o�5ٞMVJ�\���(��)C-�:�U0T�����C��ּ{I⽫�_��4�jeE4�]��լT����?Q��	�����,�A,��K��v��1�$w�mEb��I,N'������ �K�"�{n�(7)�6�˃�z�LW�� ���&�_�đI)�o�M^?���O�%y���G���7���H׻)y�EIl�^���DM$Em�"��F��-2�n.��C{��&
>�~�b+od�*n-����;"H}���ov����g�Y�o&�y6�����q^��]F�U���w����V�1-A]�����S�+��y�xQ$�o@P jȼ����Q%���u�s�?]K?�t���Wc���w��[en7+��I�_�����R�V^!�쥙~/��4��&�t�:��j����IT��FEEř�t�}��QԷ�R���"{A�j=���-.IJ������1�Xh���Ť�E�1��ts8��5B`Y��g��k�x��6����y�����a��ȿPUP~G���n, ����y�� �"���8����qY��4]��P�����1�P6+��;��wZ+�O0�����"�z������;�F	���Z~E��!4�2�� ���*���T���FB%{a���ȣ���=DE�V��K�W_�k��_�mhOt�n���Uٴ���:��%��q%����@A�UnУ�
J�LX��K(�p# ���S�b�����Yϓ,���f�R��֊�W�n��:�/ũ�dBW~����	��Xz����.C���g��=p�(1Ff�f^�ҷо�/3k�AB�md ��2�E�Qи:�1��)��f����P�����\B=<�t��D�y�m��D�ʐMh���~�]�"�#���X�_�ޙ�E��N�ܮ��8��K�,.�`�%y)�25��|��e2GM�H�mB�c�=���Ր��(�f?M�<�s=���\���aQ�[����4�����Tf2&��<f)�7U���bl��4Ѝ�����f%�s㦦AȺ�P��_�M��d�߻����fe�C �y�y�%3�阇E�ܹ��;^ vOW�n�ΝD�MŠ�y��ʈ���� ���;fD=ۺ��W�OL����6x��X����ĝ�]�=���s��R�9K�/t���B�����:5|��:,_'=���Wt�ǭo;m�CN*~�	��3��F��T<�$�gӦ�Zs�ܫƙ�r٭4������t�F�jc�#Il?�t��@�2	�O��������\8ﴮ��焯��Z |��B�$-���1*�hE�A��W#8t3��3*�BV��9�ʰ���R?W���u�I����.~�3E/t�z��m�sj����!��Ԩyq�;h�'z�� *���a�����!��~Խ�67p؋�K��������.g�{�i���;�_ɱl�
^�e�ZS�4}%���dO=2� ��~LV���V~����5
�*V��4����=�&Dl�Ww8� <Q��$NͯP]���n�>��+`�>Jz�0/;�c�Fi�=ˉ�|�:hS�k8�R퓝jU0��l�J7��j���{�x�z��� 4ݜ�z���J9�s���*�����~�.V��������!)��A�1�O)t����Y���E���L�g4c��`�g�!��Ѣ��gZ�+-��6�d2�ئP&�W���ș�R̬R�@�r7؆9eĺ�	�M&����8 t�nj�
�0K	~ڦS�ș�ӧV�� �֟�ӾMIk��}���Y(�^��G�����Kn�X6~U �o�`�V�0�R�P;�k�A�<"h-��ͫm"ٴnJ���J\/����"T"�^�&���SV���M�z��Ȳ�&љJ&�Ն� g��B80���׶Wt1�G�g�^іm�AH����ٖ�u,T`�:7J�̖8&P�K�6~��*�;{c��NP`YSǯ*}�es�	Š��Y�cA�$����9��=*��J�����O`����~Z?=�j	�-έ���F���� +�J����mm�Y��
z�gP�8��KD�p����K�di :��)�_@�3��t���g��G��_K�S��R�]S��{<��&K9��ݐE��N����4p;��xb�21��Rڐ�6�W�U���ՠ��#�3R��0\���G��-q�B�1�[&�����*İ8 ��6(�|�a������1� �N,Z��ǹ�Z�-�S��=! _�w��q���V%��O�9�
��}�p�u������&��yqhP'�N�|c'f�4�D��������#G'�_k��D��cP���; ��ԑ��0�ʕ����rm/�Y(��oefV@=�zC�.p:To�Sf'�$��{�T�P橺���V�6�D�����xF�����H �Ǚ�4j@���ȫ�l0�����PasLI\
�`eflv����<k����_
r�0�艀44�˄k�>.Ëߟ�?��dҝ� %�j�i	���NZ����w��u��/w*��a�����g�݃��>��������/�0K�~�Y�Qk�^:�n�_\3G���XS ?�$Ǘ�2�Җ����ʹ��DGr�������?r�ey-:w��Ma���q�[�_[���ɑ�^~W�,�ѻH�1;�}`@s�m���p�� �-m�t(��\?��;�에�7���Q���f>�	\w.��t}��J�=-�E�L�����a _�:��������c ��u�����$'�N[t���<���E���Ō���=��ro7F�,0Q}�|���A�������~��v�w�a'bC�g�G���cxi	�y��s� �8�w�� b�	�?6}Jz�*H������T���lD��=@�PF6�ȩ	lQ��C�K�j��-����p;�u���H�b�gL�&(=��G�����0��D�: ��q�@�����=��#��GI�8�_q�Ys.�7���RE��h���:���_¡�q�SS�3�;п��}�Z:7`3�����(cr�[�@�f��/�����v��G�s}�����h����r`�(&Q��ɱ�a��0�@ >~����Y[k�]��%��.��%���',�-��/������A\�'�_����A�bͯ��J	J��<}_x�ȸ؉11T�i	6��dӼ
+����
|/*��{���/�aϷ�tT�s��%uQ��CKe`��W�G��|~�}��L���=�ؕ�N����׻o�|@�@���J�i޷�v9�7�ԅ@O�tr;
T�>|N�LE|�x���_��C�,�v��M�gdPHR�&�r	��.�{��ز����y�N�+=�N��8���_�S�ܰIwݿ o]�N�+cb�_�3v�Kڧ~�/�1{�`��Y�Nr���.ՇE�eڱЍ"��a}7���B����LX����.RP+_H�f�������N��2 �.�3��a�Q^ϛ�ĩ;���㥷���O�lTr
���rf�y�:I�ΘcȄK�
�S~�����> ;@m�	(��bJQo����w:�S��U�f"7����M���=��nS�X{�Ӆ��>�"��/��<��Z�;�q�����(�wcP�,���Q�An���I�*�l �P	����J0��=|�$��d�h���ǾZs��UA$}�ц��-y�p��(U�;/z�!��@��G�ʵ��2���r!��p����;����;�*&�Lu��2���U_�z�7��A�v-��L؛�6׀~}�*�3��AJ��,Ԋ�s*��c�AuN�f�����۸P՚
jc�j�3/�ʄ���I)�`�u�t�����"f/���2�D���8 N�������j`�r���Z�t���F��g�Kb�m fRϵiJ�!̎���~�p�7|-�M��b��L.�Fj���^�6uI��Zf�[�ָX���@�^Z���<}�U�Z�˪M�@#)8݆�8k���,��Y�|GNO1V`�]M�2�Db�ૺ`}�>hx��>k�Ʊt�-IC�Gq�N�$Г�Tgi'��a���� c�I/T���/���x��6��� �٩����m�BR�>�(3	��5���$�^6���w��D�ۑ'�0�����
�pERPyL�(�D�65���/C�$�j�
0���J)����߂�E־}y�R�,�KJiٿN�d�g���y��s�-!�����^}���r��`�[�1�e/���-��7VX��0v�{u9o��?z�?���8ٵYa�ͨf���p����ӆ�l~�(gmI�<��>��;
��+P�i���a44�,���U����Z�62Pu<1�|�i��-�;�/��R�@w���4�w��9^9�M���B�2�s��
�e 7Q��Q�U)w��� pF�`�����]�Z����� &4�ŗi�l��+K�F~�{y��C�-v��y̅iMx_�k+��BF�u�<�q�w.��o�=�@�U��갾Q�W�Q�8�2��7�g}���$�.R����U�����@$O��Z=mt^u�V��/o���+x�l"լ�wI3_�[�Wԣ�/���+_5}�D��C�$����▿��Of�(�u`#n�O��9��W���g4�)��2N���{*������X�J:�����(�d;�J����'^;z�K�1�~�� �Č��	��r2�' 4�c�$q(����#�^n���%�Bhjن�>�ϸW#��"i��c��������5J�kJ�5�(y�6-�f݃�W�cb���&��G��J�m�Gu�)����V߻:�=���v�%��#��6�KhK	� �C�u��85��u���{	_���ɨ���H�^�&]W�/�-=ŧҤ[l�f�:�i�N-f��GA~q�u����7�]i��I�*�K��M~q�^#5�t�������	�y5z �@� ���t)(�c�ێ���j�J�P�����oB[d#8LׯH�⻼�8{�I���yl��2˒��%E&�o�oK��t��ޮ~X�_z�8�|�d�6�Í��PW��1\��h�۵�漦���\�)����w�_�c�"���B�va:�� �2�W���';	�~͟����
5RE�dJ�����ZK+��`41EC�%ߺ��k_���^��1�D����!�G5�͑'`hs炠3�y�+l8۱��������[�/[v<�!k��Y���T9K�k���'Ǆ�x��J�d�8I$�NU�QA؇Jd��6�:6�����(�l���}��n�W�l�JVOݫS�n�Q8L�K�&ĔA{����|A��
�>k6�VLNq���*����x�#���b@9���*����i2������<}�mF�ة����U�'I��#+{�L�P4}�+�������268�)3��:(�-!U��^]RcC1�F��lƒu�$��N��A]�������D���W������S���BMw�/1��I�I�'h$�|:鏁�����G�[������@�O��~δ �Ҫ!g� �4�Q���~F��/��E�\�'�W�),���J�2�u|�Q�j<�����͜9:L7�)U��	����5��/��}�ⰾN���UL,u#�'n�g��g�[x�o�ˇg�m:�OPq��Ԗj�DY�����ӡ���� :�����q��
�r���0���[NP`�������"~J.w���)>�~�XpHeZI%Q>�F�%����~N��f�hx��S	��a��[��|0ܦ��0�|���c�1*B�?�XJS��,�/FJ��Q.bp��$�8=���h��i�oD�σ�$U�.  �W���b�� ��FZ��O�9�=
�sʸt{A�'	fy����O�����a;�&bX�{�-��~�#({e8̃J�!�r�P6;�@���aiQƜ�FxT�����v �dw N�}a�3�6���^����
���%���tM�8�6��b$  �I�V�9 �F%X@��E3�%������]�DY��J+T������S��_Q��1l]L�e���;�
Eנ���kDFj��d�/Ϡ��@��Ρ!!�n>_���	�r��5]�H��\�b�|�̢(�0X�S�s���F$�`2����{Jk�ʁ[6��V�zH�y�=��QP�!
� ɻ*��gb�-����-}�?�DGX�oc��
��F��P�W�o�h7�m	�e,�b�k��Ą�h<%�������ʶ�<Q`���Z"/�Տg�0^�{���a�s%���l�������Q�P�"�ߛ�R�
�լm��"y9A=�@xb��
�;ٶ��#�y��,?�r���lBS��f��9J;��.�k�埰_�yf��\��4�g=s%���
,�D�ԻJ���d��m�1N��k����k������;��~"��6��l��iD�}!�qE�����S��5�����V���ب�A��%���e񺯊�YK>��N����D�����B��(�14X���Y�i6����F��s%{.3ᚏ��������0�f�+0�~���:�9����D��\�#�R�?w,�j��l�P�/l����|� cA'ЦG�{U��X�Z!&=�^���\�,�WH�Ls;9��w�Dn��sC\��LH���Bw��T��5��H�4�J���r�+x*ܬ#dl�,�S�k!���_a��O��5�S�"}���vL�	r��ï�R�������P�ǳ���"�E�{��i0�A��=��`����U�59KT+�H� ��0Uf.��#3	�����]��F���P8���/��{����%���fC�ei�}ɾ�]c�¨�-%*#�d#!	E�6#K��}_~����^��ԕ�>���k��y�i,l�E��p�h�:�Qe5��4�Ԋ?ߞ�mw*�t����mM���DYfg_���d����O�u.�J���'r������bA�A�js���� �Ӏh5�SC+���ʟ���8���Φƫi>H�@1ʽ"Q|����k,,�`�$�� *�ߒ]i�ʿ�~J���S�м3 �YF�+'�����`RE����>���H�f��B� p�;��Bo�vwQ��K-x���92w6�Q �,P��u���K��A����i�)!��C�3!�:��+��nԠ���n��ݷ�?9�-!��;43m�s�V�.V�AJ�;�"����]������'��� ���n�*��#�S�M�@��Op�Kp@�ټg���nnZ�w���/���3xV,x�fyl�-��R�����L�$P.�*s;�{s�(�s_@o�b�����&\����}ޠj	{Z׿�ê�.`��w7��{l.��ć�,C��O��c"}80�aնH�@_���xm�A���|o;$Q���r�R����'�
��N���sq8I~p�P6I��,@D����7;)�^���r��u��y��Yz����Yi�awO=D�P0}\/G稙AV��VS[����n��J���]�*KMBI��9��LJ8]���<��31��CN��N<
�+@���Dۄ�|��+��m��7+���W$s��W�5WQ^�ʹ���A��7\���Hh���f�d��^V�qm��^~ {}����T�+jmQ�<��'����� W;^�	Oɾ�u���jw�m���1�p�!�+��#���Ns��'��;z�s���������%���K'��{zz S��P�K���"�7�i��q�ҽn�8%�7A:��M�j��!�:�;��*��e!SU�	\��o�9f���)���u�c��R�#3�oF� �8������@G���-�ꑀ(M.f����3$UB%!Y�C��|Dn�	f��j˭���왯�6��a��7L�DlAy^ڿr%�\.����|?���Jc��M<%^�m�^�ؼ
 �4)�a݂�FN}N����a��f�9h+=�ҕ�(��R��|>�*S����ࣰ�\�O�{W� j!� D��������]���SBJ���,?G�܄���'�ɒ�ơ+��ӫ�n2��������"獀�����ujN��>�ۍ�X�4�.To�м��r&�M��їV��*tQ���@�e$k�2��Ea�j
P�q��y_����X�{-f0��c�����x	��ᖼ�eEM�BJg��!���֗i�� �~�$�R;���=����'?���
�>�����|�j�Z��.Q�D��R}Z�͖'?��>�,e��&
�+˛v���)n]�]-�����D$'z���y?<_x��C�X��]HyEj�2�,�`6�7��mM�����d��
�e�4���ܦG�o
�=x��r�	��TN������#��@=�r]L�>/���X��隇���,�QdzUϸ��e��@ ���������u!��h]�0���"��	J�zru�^:)J����|�f4�g���ɺ��W��,`�⽻Pc��NA=1��ح�����'g�O�@r�T��?���F�?�~�@�b�=�T�6DKL~�Y������5��� �F�ų'�e���ϟ!F�=�T���P�:���{"��|̃i>j�Rb��m�}Qjʗͫ�P �
�J ��v0��2r���;��r[bZ�@�e��ua�.�ToQ���D�l�Őc0t����jPҋ���&�d���!�H9he/��`f�s��>�8�/�,��?m�FhO��D	��v�����dʔyv�/�X��La��k���_K$�RV��x�IYEW_u���.[Z���Q�3^R�$��]=�=�҃`?���̾��3G���P�;/��f�(fiN�?SW�%N �j�����^�d_�5F�1�Rs G���S����9>����,���y<S�QKՋ��yM�FMsy�;'��#]3�7;{�u]�:��3_H��'%�k�\�t9�����RF {Ӹ#P. �xx�n��Y�e�
�~�,F:"LQJtCG���������ј��D!i�ٞ���:�&�܉.}!�w�>�>���.cn���ׁK����_O�l��o7���X*���8��%���mW��,� s�.��<�n\r%Jϯ�"�hJBQY�l�B
���t���)8V���f���ḻ���{���C{UlMG�M�i���}G�y�)��0�a1U�Y+�ޠ1�б�RA�fd��i8�G��1䘃��7w��i9j�dQ6��aє۟��N;v��?���Fy7�	���Ʒ���E�;v�z�����;n������x�K����--d��	,~��,�g���/�%TO�&9��oe��G�I�i7n.�p�wd��AJq!3���S�6tU�M���hzb����azQ� �7'$���r��qE��џ�����},�e���[�t?# ���W^QS�s:yV)������l��S�Y&��^�Z�7�hXIY�X��u�"��J�P_
n����#�x���'��sTr+������8HE�9�|�5b��$@8/er1c��(��|�qIk���ZW���J�$O�h懓�8iYI��+,m���o�/N�@$u{)��X(�p�b]Z�CG�cs�m��J.[Bx�?��"ק@1����KԈv(���XQ�P�^�W��ϻ��5(��B�Y����i$���E0�����g�*<�EVY�Wϳ�sS�_��3::zT�^#�ǦɅb�;�QjX��%���Qa�D���G���cJ�TF�^���d:�I��P�>�u��̈��U�@��p�෼G�ۅ�P����x��z?�9�2-���T����G�
���b��ʖ��B�k���v����}�@|<Aj|��	��N�s�r+�1z'a���"���m�m���"Z}�&;R ^�� ���B��Š"�s<[�tb��^�B� �>^)=�C䝛� s��p�2Rͫ�i�BT]���xux<HP50�ve�q�%mM[�W�^�Sٽ���h��E	Q�Ά_�ۛ�쫺��L�$�Oz�a��]�y�OInM���L��:{�*7��Ř�㣡0@�����R� a�8�:����])����"YV�f�Q:)0�!����OC;�dG�\J:+U�q�����(�[e���ӣv�!RS[�~��l�K��/$�u�����$$^��(�$�vx����♸�>L��:;��5��p���>����Dw{�I�  aW�e\q��xa+�O�?DKЖ[��l�������-����3�u4��)%��ב-[>�Ŀ��լ���x@6YmM^�fg����ϥ�����_K��d�ypZ�Dqril����j�Q�B��ӊ_��/�typ �2���Ж:�a�:�'0�N}��D�$����c�=�����b����D�6m�Mhj���Y(Q���p�)P }±�7�u�ӗ�5�5�*���X��a�x��h�ۯ�_���%C�Pt����`�"�:E�Ly�跂��"S^�s����͗�	�X�#9H�w(E���ZJ"r�"�F��:�pV=���n
"ݬjN��w���T#��6�8��ٰ��G�K!j��17]�9:�Z�
4��׮��Te�9��������wfbS���J��Xi��'�&n������֗�B�?�ٵ��J�N�'��� pv�j>��̸"��Y
gu��<�R�Ͳ6L('��a��%Y���T9���p�ҦH�O�e=�R�aQq�v�"Za�
���3�m嶘�A��k\��0eO�]b�NÔ���:vh?�e+Υ��i���|M>Ӈ��c��Ē��t�����>�,��q��ocϡ0��[������_��R������,�uf�pַ��|:A0��CA>����Vx�maz�	��x�MD�*H�p>�/����}V�٦X��\�VU����(FcVr�l2nK��@`?n�з6�r�4.d���%�j:�%tR�*ƥ~V�S��D+9�}���g0����{Z�6`�
u��BI<������EÛ��hnR2n�����8�&/C�b�H�(�Q�-����oiM�%T�ky=ۮq��(v@.^Ӥ�:}y �V��.?1���� 9���y�<'X������>���Ÿ��W%��h+�oj��2���ZC�N1[��2���¬� Lልo�U~�c7�h&�o�����B���L,��ن��ٺ���EZ�r�&�;$_��o�2�x�"����y�#�'�mRu�֎懎�@1�𙔺i�On�\�0{���LE/MݯHЍWc�K��
BZ�p���ᏼL���gwt�7��`
��;i��fώ�k��O�jbY
����-Yv�1$Yܐb2�
$H�4~��!O\^7������<ֽ�F�3am�K� D����>�;�ZPm���3�kotE�})>mQ�4nycn$�Q�vU(wh����VAg���?�1OJc
�A�=H;@�u��X�������=��SE�q�Iiۓ;���!�r�*��Ƴ�GM�����ulp�	 	_�4�(R6��(��ǎd@�����mb�U.|5�
mO��󖦚��J"ذ8F 2��z 1�b/b�ŧ���O?z�$$�Us�&{��}�B���ޭ�i\-�5a��s���)D�a���8��!��z��-K�<��-�W��#/�G\#oTbY�����F@��ý�w�8](��7�J0K�ݪ�w��3'{�)ϻ�`�K~��z�Qw��/�� �R4a�駜K{��5r��vM! Z+�p�������ӈM��*=�4�����&�O���:����?��{�������3��<V�Y	�����]Pi�����4�U�Ƈ�LZVtitF�XQ�d�x�`�
��)��<��z�	M�]E��� ��K�"�yA͠s�z����:�b̰���I�i��w�,�dU��j��F�Ϊ��`n7o��^��5�qO� I{��j�i<�F|��@�j{���o�Z_��d�H�Ķ�Y��������k\x�w����K��d�>+���.��vHz]�:�vO�B�H�2����S=*	�T0��3-u�v'����7n�qwY����$ z�ޫg�һ�ݨ)P�;���W�n ir��<u��kT�+��d!�b?<o�`ꗱ�T�p��{���|������E���oL��k��9�-o�hStyeA���LtƦ�P�j}��!/ͺ$-q_��c�IH�C`��i������	�)���iY�f%�����zfQ�F|Y��\FE`�[*��"�E�.�èB�g�2��b���'���cG���`��QBp��mH��>U��2Xp��ǯN�P��n#k��y �d[�3-�iJ:��"Y�4���˂a������g��=����*R����yr]���*Yy`�<`�`7{�� /Hy\�a�Ɵj�Ú�}ָ:Pt)��,�=��L�
?����z,y��gf�~�D5��oofy+1�3�yMӡ���%�Xn�z��ʚ��ˮbh���b�O3h��%^�Sq��	a ��=7(�x&6A�lT5���ٽI��ZBV���H�jͣ�Y�>��AQ \y�P�]���3S�������]��w�R�e�J��A����V?�:�5�rZ����|e�[lk[���q��iGܘ��'��;���2"���P��1����3ĳ@�>��k�,�\��pEk��ф�x q�4NKL��q�/�0)Ց��"�)������/�$�Y�ƴ^=A��z��U���z�}~�q]̡U��d�Y?�)��Hߺ���y({�8��n揤:�tB�_�(�L4$��<�O}�E��{mﯰ��`�y�vv��_Sϖ�`��1>[Z X����\�H�|,��k�'��y���!�6Jv�;�j�l�s-�7KI�XFv�
�u����h9���X�>�+Ϳ'@u�ɢ�UQ���Լ�[�H����#���J_
G�=�DH�]���i#,��k��q�h����gP��I�:��A�62<��&7���BI�Y���A�Vt�P#����bo6�	n�� 4��Q��B&��&������EK="2�W,�~N{����m�A�)R�����0��?�bM�@�|�2h0�o��\�ȑ�A6@oO�`����^��}�����u���w3�x4-b07��Ӝ���e#'�T��gu �*����Zg�_���O~ڐg�j��<�x�q�Ao�����y�j?0���Y�z+�{)8��,��x>(L ��@f>� �:qI./��q�a{�l�>D�:��O#T�P�df�nC�r�]��gI@�&NMv�@�F"q�F ��7~z�i�ɟ`P� �v�n�w;T���)�N�y����#-G��E`�o�+�` ̟�>{4����>�H9l]�A�C�l�&0���Wn�a��'�+�^��iG����F_�g'3����p0�v���j{�f���Q��I�P�i��*HxՒ��hc*����~b+��Q��P~�T���W�&��H`v�4VR7kuҨ`
��{����_gP����&�s��E�}>O=yȲH�4,=�@Q��O�f���������oщ��*#3a�{n�=�sh!;�x��_�C�"*�Ť,�w(Z�T�;�	�2�����oB��#,J��h57��֋�$?:=�F���y0��/T����l�D���"J���67�Hu�[�@�7Q���7��+i(��;r������W�;\4Ү?����CJ��)����jL^+#�v[C�Pfl2��5Pi>,/>�_���B ���R~۾B�p壻��iӸ��5����PR+kQS�n��/Fn�B����1}:��ӈ u/9�K}��?�L*�IB���Uw��Go$��^���̽#�0�ϒ���_l%�#A�g����E�:XaЀ�}��������k�g�r�Kg�VG��5|m�2x!��5��OR�=md:��{���%~�dkH��	�#��[���r�_�ڄD?����l�( 5p.$?�*9ѻ��Ч��Z�����>��veϋb�\v]0[����V��Í�5���=�20�bI13����=B��v�$ߡz������X��ca>���
�Pd?�N�3�u]�s���H�xZSo!��=g�vstz��E�����`�Am��@z3{GE���%h�FM���w�3��+�$<���{�:B���_���@ӡ����U#鏲�3�V�Ԕ�����2�&�r�&7����ѐ���3D}�}!*K[���Kʧ��#�m{6���7��3O�Z��kr��gO{���Q��, 
��y:�7P��Pc�+����45~p����mp�dme�5%[Ce�E�d �gbRa\U}D��bTN�j����R������8|������w�8�j�<[-ǹc7BYO��\�����A>��Z������k�f�\� �I2X���y��.w|�)<��S�������
��!0�E�������R�_��|�W'��� H�2��po�(��x]#/UFʩ��V�̹�"���^�+ Qn���>��{����R�)%�7�֯+X�#��Z0T�U��Y�}�S�"D��a��^$�k�E4�v��~g�у�bS��1���RL�Y��g�ٻ삉wv�0���<m����4�/K�9���J��R�8��94)����Ũ�cu{��~�ә��3���;s��\�%�^L�� ��bWP5��u�Fz
�ǒ�j`�d5U{�F�����O�zg����&�`�9�p�e���j�d�Z���1�cfӟ��p�o�2�>���)i�_�x���X� � ���$uzc\�)!9/F;�jEgqa��@3|�&x9Tvn��f�w�i���	�l����Ҟ�0�Oj���y�M��q���@����I�m~w���Ց'X=Ýf����Z����7�=,��tMѤ�C 9��5%�c���un�)�Fw��}>�����܆��w>���	�8Rd����d��Chq�<~Á@%�<<t��DX<�HI�#���5�>��$.��<ñx�[��龍l�Co:%���*���$ HF���?��Yޕ��K�����x��:L.����ЄL&��7�:�Of%�fM��2rT��@n��)���0
�Tm�����sj�����[#���26�����e�l��q�.G�e�Bȳb$��'
��Nу��n1i���ֺj.���X��$�� ��nsk6L�2��_� 8_h� ���:Y)v@��s��x�JX+ʳo111�v�^�@%�*5���3���p�c��_c���\W��5 qu��s~���'5�e�"��8Π�[�$9��/v�ߠ�ђpw$��H,Ҩ?�Q����ɺ+�>s} ƍ*��E���0ﱈVo�P5Hg���s�:��A�]�:���+f�gg�E�6/G���_��m9!EE�#��/"is^�{�sѶU��e��E��*G7��)`�@EձI�I&M9�(7OF2F�]̣������X�>���c�˾.<Q�[�L),�?d2{�isc��!������*�16�]k�P���̠�cpaq�hƟ6�jb�T���T �fy����f�Pԥ'?�~`nu����%�4��#&>������ЋP�u��X�M*qN�!q>���`��)�ښM��gE���Jg�m�ͫ%i'��p}����:knV��bO��Em%[��4n�+a����>=���H�nKG7�ڪL�h�C�5��o1���b�n�ׂ��TU�=��������(��
��%+�i+&��7��h�a�H�0k潻J{=='�[E7ި
�[X\W���.ǯ|�Ak
�Ǚ��4��������*@ӷ�$%G�$�b�ڜR�t��{�ڄ'
���!�W-@�O��S{���~Ku)D}�-;k�*�m�����Ru3BU�t�c��i���>��U�RCk���h6�w�;|[<�L˾a~sYJ$��P���6��բ�`}x�fS�V�y�Fk�`7+N�g������BN)r�p*� a�{D�����o@�]�172��#�5����z��#yy0U�C��vZ�c�,��*�є�l�ە���n�&�F^�_Zpc�G5�����^	���Y���ɫ�r����FX�)уg��b�ŅL�&r� ������D��H��
�O�H|�e5����WY��T�N�4�ą[a;����?������yE�1��H�Fצ�r���M KA��i˄Ռ\ڕ�Q6j���YR�Y�19��K���hf�b�NYm�Q��/-�����<�C:�iJ\�[H��FB��/�˓��4�����Z����bIQ����eY�Y嬀��<�Kk2 <`*���W�4����l��}~L�K�_Ɠ
]�v���of�#����C�P;5ۂ������u6�!>�?�(ٔ��>w����M��+b����V.�HJۮ��@5q����]�	��qǸ!P��P���[w��� 
��Y�F/�ا�����Z�>��_w���oi#��<{G��&��1)���u��]B�m��	ּ7#A*�-X�U7���V�9u5��y(4v�ă�C��v�\�,Ԕ� �c�W%c���
�-���Љ�3O����Z�|���v��fo.�����>�M�x���&�[y��f��S�M��.�����ZQқ���#5ɹ�Q.����-[��� a��Q��5��#�#@_��O��,=d�j=��'��oƺ��Q/\j�O� �{"�D�2����/��׃-�����Vb�7�pV�fv"
�-�ܑ�[���ZS��jҷ</7wGñ��2�Z_ RbN����cK-��t,-*�) �ӻg��jMv}R���J^=�]�ɔ8Z�d�
����\��R*�Z"7U+B���If�U�f�{c�C�{����Q���@��;��
T2�l���*T��]��a���ތ������JᑬPB@v�z2f�¼̆�R�м��V�}L��q�5��ٺ�F����<,[���E�=��	n�"ˡ"�������( �K��G��C�幥��m����"�����9!��|1ȑYf#��Li���*��<6�V��H}�Hӻ6mj-�§��jBl9�Yԉ��k8ܡ��ы4Us<_v�%đI���R�����AG��-LAY��V��zŭ�3\����þ�m$��{�����z�e:#�+4v�~��[�m��!��;'9� zp�΃����#;�e��U���c��uP��g	�LC5Q�-��]��jp�Wvg�I�U�9u��ï��z+5k�ut����1uu�půs2��^����DX��aUڼ�ld�鬧WҨaE �G��x��������TQ��1F��{H"���4���+�o�P�������/!�'�o-�Q�
M�FT~�}�y��sU���8��(f��`�."a[�t[j��������T5w8+i�U��]{4��Y��ƾ_vi���? z�u���׶��_���M�ҋE0��x�oN�/��>�� 7:����� ���׈p=l�����΀*g[+��(μ�.���7�:�N�s��}�����V�A\�֓��jd�pgVV�����a����=JCs��Q�sf0��Q��#Ì�?~%���+���3;���}<�����tM�cy����A<$	_��xgu�z�^�*TPϲ�Ok��&�l���>ͷQH���Y?�d��v�}r3܍Bh�>
��+i�/&��	��Z�<��\�?w�X]t([�8��`����Qlf�)�f�3�B��#ic������n�on�(7g�*�G;?<�whqGJ$Ǫ�qY
���<����N��)G��{׼{~D'+W�΀��
��󀟆ktu5im%��Wb�]-�۬�֟?��/%֓����Ê	� ���7���i���2�u�[P����j%Q5&;�J5�HJ�-<�a�|����'5��cr-]Gz�B�X����hX��!�A�7�%��H�J֥���c'p
����Tpb���M_�[!h`5�O�f�MF�]t����|���]���ӳ��c�K���z�^�~w�I'��K���c����J��):������Xz�	�����6!�?�M��6t�w��-3��I!v~�v2�s!x�/�+2�����3�g��i���%��;���W��"/ !Ժ����3Z\W�E g�w;6��bJƖ���O0q��T�jo/�!������Hn�j�+���/�V��k$���f��y ����<Kq�Y��.�j"����t��L2���4+S��|=jo������D���?t��N]?�V tZ���n���Y�&<\�|��'j�����4YYh�(|�3� x$��P�����
1J�x����qJ�FN�fH���rt�@�\>di+�A=�G�Z�_�x�_�UM���/��QI�� �;,�UVn�Jc?�l0/{�r��Y8kx�mt�Z�6�)�>�z��+H��M��S���}=sŲ�,]>�m�kkk��`��VW��y�Q��1��6��H"���	W/��hn6��ΐͥ�
|�.��,|�\K��z?���b���8W�ҶPp��U�������RH��\2�b'�����Wj���*�Ԉ`��Sx��������f��(.k��yb.d��尮��6�q*�,�yK�_HM;��K�qo�sߵ#��@��R�M#��Q�?�uҨ�����ed�Z��C���p�aYA{�m9��B�F�Q}����o�hը����'�����>�	��1�٥�JC�cXQۚ0��ѻ���x��T\�H�� oX��N����S��?%��UT*�㭕#�q�����jꜬ>n5��mO����Y5L�v�@êjj?&V�|ˬ�[�������1U.��q0�O~�Sᡭ��z<n�����`"�����t���gЈ����Ua!|�x^��7i����8>�,����y�vA9P@�z�׬$�j*�
��D�H�����&�~�l�|V��@�~㿄�[�`��O<�(�d�߲�Dv]F��P
��B��7�zX�,������a1K`
_�����4�u���N���ԝc���K}�,r���~u���p��,�}�e ��o]85;�Ĕ�"�@�K��bK�ɡ�죸�e���N�|�J�3n��r�`R�صnmc�iW688t�kCOO=[�u�2��p�x�K�؇��|\62Yl�O���0����]�fjʯ��󦿘`hX�~��G�p5�i4�]=�:��
������:F�^?�fNn�t�pIG"ǹ�>,vo����a��?>�[����5�PJ��Ћ\}S�����	FE��cZ�s�[(b:-lG��]�艠#��/񷜁9tX`,��?���>�4�i%Y� h> 1ZY��B1Mݥ��R��v:�8SR��F��Y�~0���mۨ`@>Z�ٙ�s�<񭭩�?�J��m� ���gve{]���i��ͼ߻������q)V�5�A���#l�}s��"�W�`��s��,l�;�c ����]�kdK�k�ǎ�.!�;���\�hX�8�/��6^^
�eg瞮�2���S���c�E�s��JM�KAHX��߰αc�ﾵ�{۴�&�jc��b]�Kɤ��9k�R>�$�k#���+����#M LJ�����ƞ����V8tc���A͖�>t�h����#Y����k�xl����v�w�����Y����ް��s����;��R��'[��䥜�k��X���/��r�]�ģ������^���`)�	�VA��Yֲ��׳
�߭z}��}/�bh��W�,y����VS��k�eD�����o�7[/,	A��n3�NO�9��ïBWy����G����Ѧ0<s��(P��Hp3��X�\��`�L���A��J����`%%H��-����|���]��[�粨ۃ��vL�<�1Ʒ�L�6��?̵W,��I)H�\7���<_���0\üԥ��ɝ�k�S�E�.p_۹V�t�C�΍}��#WC;��']W/pN�5 ��#�Շ&��cgd���`�7n��4�����4���>�
��i����v�y�<�]E�y�^�x���B��~���GT>k�cV�06�~j�s���ŴlP>�Ý;[Ŋ,��"�C�g�.{�~\ы�(�%01ݥ�T7���������ū+s�g��p,b�rҠ�����_	QF�{�1���&n��6�I1¸b��������, �f0��S�_S�&�:�1�;VwP��^�@�ha��C�q	9���t�������F�&���},��u�C�n²�R�t��OPY�U�U���K��;v�?TM2����y�Pw}������-������,¹	v�rɫ��)�@����K���^��i3Z��A��v3ͭ��}�C�o���k���k���4X���뫮#'���1W�5�x6�� ��ܼ�����˓m�e�PF�����z��ʍ$��7��KJ>-#��=��i�K�5���ԡ� `n��K���k��B7�K�KK0���b}��T}\��7�6��-c���pw���e�� �?Z<����5Pn#~|����vM~݌��gS�`�Y�8��\Mn�=gZ�aչ�RZV�T�D�#������7�x�0�F��wv���N}N|\�t�י)�o�w�9��cc�I�_���c���_���x��8u��6������^�S�98�"D�nQm�E:\���{i��|��O�^g�~)J�S��r�K!�=���S��m�K�8?[�G�/��:�E��`>����>0�� ~��A���L˟��T�>:#lI��D��l��ͺ�1��諔#e7F~<>Gx�-#~�Rד'4�R�:4F���̓�Ca�;C�^�~E<�2m1�����h'�Ӯ�T�o<�Ɠ�[�D?0`SU��Y�n�Qz~?���4c+*ԡ���A�ǃ�h�Ɠ������}�q�hR0t/%�!�������i@ּ�>;��}��V7+	��ƚ������w<,�����Kg64�a�`R��Y{S�������wR�'+�[�'�`��et��*-̍�咱�����?��D^�(V���v��3H�z��2�T8Rs|��"�:���ˁ�kg?�D����?����{���O�X�#89�M��Ժ��WU�G���T8��� <�+�,X�'��ݮ�[�+r�K�A|�N�>y �U{χ�Z��_�2�h���k0��O���/<aDS�U���������Z�lJ��ol͏�m�U���V��Vmɳ;�����pA��m��P�/j@:_�'so��g���54��H�ռ�F���nJ��<wO_�/Vgˠ�a��.��J�[2�ZY�l-�h ��
���V�
�32���T��$��M�w�G�`�z   �ݭ���f�7��&�qz���r��/6���я:򃞃�hk��g����NNm;J時�Nt��Rn����Ϳ�*�"7���"�"N�0��s�,�LG��V���/-ۨ&�'~>�;����R�Q��H{bIN���� �mG�f���*[�R�5�Z���K��i��!z��b+e��;o��x������$$��0�)t^���4��_��+-[z�5��VS�wW��ʑ���x]�;��2�@L�D�?R�����*e|yrg\E)�x��)��DV����������bP�p1�����U0�N�����q�̕���ʷ���0��G���F"Q��^7�a0�^@t���%��[�ԽN�<s��	kߨ�j�J���dM�S�����d"9�����Y*n m������l���Gg/��mZ�f�6|����N�p)hƥ���z���+V��~s�t�	02��h����FX(gŗ[��Ġ�Z����Ɇ���F�(+�H������I���/��e;JԘ�V}T�q{���(��e�g~\BO�6����(:�n�k6��e���99��}��.���Ҥ�%��[1�jo8 s�	�����f�ry-t'=P�H0����H��9u�,��IH��F��tcN�?j����*�������S��-��'�����3x~~~���у�(�8��0���z��;p�k)����D%}y�����}\}���T��E���h��#:�A��r�����UN��[R�}�x{�=���,,~N�@
�S�iwZX"�?][��$�u���ꕘ���u{�y��{��|N���X����qm}��Y7+r�UQ��QjX8�՘��{���5;6�`\�B#�`��T9$]�O��Q�LB�ԩ�T]x01>�vR@����UyI��P��O���o�
.�k�P4�}�E�eW��̬���77����wO��UG���h-�oW��X%�L��!P����{�5�^w庻%{;=���|}MF��7WLJ���:cW�|X�8����w�糪���]r���;��6�Ѽl)"o���,.Vy��P�z� I�2Q�E|aJ��rh�jGW�A�&q��.ǈ%��T�P��.�|x�g=%������^ڒ����lQ� O��m���%P҄,����||�XG�w8����<��\[��۲4-f��<���@�>��c��Ѷ�C#*t��$�O�w�6��]��K�ђ�s~�fW;q)3��>�C�Y�����A-�Ǜ�S��>V����j�9���
#N����&�d�n_�7��6|�$��;��*ka<�/� �g�D���ڏb�\�/`u�v>�O�15�����k��;v%� �c���{d�d�9���c�_H��6Qp�\���p��kx>X���5G�k4Nm�P`�E�Tt8�^��O|���ީE-,:<gHB�'5��Q$I�I��6&��O{��ׁK;0��$�ޒ��!�;�(�^kZ����Ky�Z��N�jhOn���J\�G0�!O5�����y!��������E�ꀢwS���&�o�>̓�17�l�_�[�](�
�"_�ʢ>��cϊ�C��À!�	zy��8c{\�"Y�,���#"����o���}�֒��+t%��H��o�4(��?K~G
��-@�?��rG�Z����P4=�'��ܰ ��û���`��Kp&�2Z�T����X*��-v����=-��
���g�'������䨰lה�)]�MN�K�"��A[�{��.�|����4C����b���%JTY[[j�>��S-�Z[�>V�b�18�=w6QA	,`?:�f�֯pm���#�+�.�FO7�Y����T�V��O����r�l���Ӱ��2�$l��.Շng�]|�z\�W�2K��?1=�[�BK���������:�quq�c6���ʨ��IByyC�wq���z@�wp�/ZIi��N���:���.SUE��Q?w��5:��\�����;Hh8:܃�HPsE	�o����]���_]}���I(��*J%��5P�ꕾ�:kk��JsZL�l��y�4WS,N��66p	��
MO�y�L�� ˶x��~=:�5:ܴ��h�vw�
��u��W�X�T��V����u@�W)��/=k��N�����TR:虓�P�i9������|�/�ˠ}�7�Ι��U`�1�&�����b�h{B����Q論�_��=q5�����Gj���*V�;e��ȹ��Ζ��dkZQx�oҴg����M�>������+� k�v��њ0cK����*�x������ǆ��{wq��w��s��4�ͥN��pxe��w8�k?������@�{ۓ	g4˻`�s(Ԇ@sҘ�\����l�>`0Z1x��������b]i��۴^�'����it�jV��\�rs`��\�Bu���m�	mL��f*��=7���[5s��]۵����i��������.q��)�ˎz(<��`h���P��O�o�s��'Iʰ�����w�ؽ���x@�ۤ�O�>ͷ\���wc ��2ld��?��S�˖�1 �?��W|��j�|h�m��^>.NʊU��W�0�v�ua�p���X忨�A�U��^c%�[��&�߅z1���xJ��9Ƹ�y�����RCS̴���V �߷����2��k�� e�tW���MgU�~�!Ei%��E���A��[���A�[$�F����F����=���χ��쳯k���{�;߫,�2����H۝5��7Z��Y�VF7��^�k���+�B��x҆O�R���LWr����IG���;,�Ŝ(�?,�Ṉ��~ޖbtr�}��󇏱��=�
{�ҲC y�Y���a�Kt�[��@?O^>$��x��\��V�����7���=ϳ���*�W@|H��zz'Wm��4��P������܌��|�Pd:a~�]v��M�VI��$���^s�i�X"58��xzz� M�	�����=�v�=��n?~�����C���q��/=�K_O����hr�s��}�B������U���59攢򭖓7��mc�f�m4L^j�-����j�jJ�8o}=1� ��wv6�g��c��G��|�e]��SD1H��y��V�H/x�bDc��t]ʿ3i5��vC���&T�y�C��5N �)��QI
��C���DY����@�o3ޥi�$�/^���4����z1@��V2���jb���i���������i�/��ތִ��̧�s��ܾJ��#,
�I��n�9�����2 ]ѿ�Ж�߈����G.��x&�j������ROk���6ZVx�#�=� 7�:�&�*Z���)U���R��Lmd�]9ڢϑ��d�X?�z�e5��-����	��E�iY�z�����s��q�>ŬvY722G���k�+ú����:F�:�pd��p|����Aj;,���m�ڇ.g5�Jļ&K��0���v��H���V@5��T�J%B�"u������golile%'���ϥp�7��s���=��iY��8����#�p:���L"_�=C���s�^Q_�.�;~D�!�|LY���n��U�&�
�a�1��6��!]�ߙ/]'��hS�����������_Dy�5P`�j`����N�8X�UM�z"�{U�5�p�,8�.I�L��_���߿��q�Ve�EO�O�KT��&W��������x��'%�����K&���	�o��D��%k�>8v3@�pU�l��d�
L�LGߏsJ�k���<c��R���z�4����l����k�=O˟��.u��|�8|l_ڈӯ�bp����J����ݿ[�ؙ��ݥg��"+tm��k�m��A3��]l3��~.�����~~v�S,���~�8u�;\O�j��X?�	W�5$���o��S���~�V�����ݲ�m�2B���d.56iG�m�\e<�D/ � ?@v��
���K��g�E���R��i�}p���0}�7/�O�g�N�$���5�����Q���H��ʩ����_� |�]"NQ@�1�!y7�n�ka߀7�KN;��1-�G8Gd����!��罓���,�����\��X�br�#��!�N1�h��\�m��q'��&�A����g. ��LF2b%�%3_�F{�F��a�����v&� �V�tU���I��F�fy��6z�L���(���og��lZ��AC��0C��0�+�ZN�~�s�¬s=�_w��pR֕�d>S�t���nS�����}��`����4Q� vN�6\��.��"$VւcU	ls~�^��Ĩ�l�F����	�����C���y�s�?c��v�߯=����,+��s޴�<4~��N��B���iF������+S슊}���1�gנ�� e�UWg?���.r؎�-��������aݏ�$��wD�{z�+�:�+��d	���G����p�`�"ȼ���P���ʭ��䎳���AhX�o���kŻ:7�(��I�<H8��	�@;��w�`D�	y�i�Z�F2{ڤ�tv�O�Q��o��p3�Ou4c�w����1h��m%�k���������㜇�LbD�eC�����ȶ�b���XIp���������9Ek�߂Q%�����u�1V�}�����A�">Ԋ��]�l�G"�Ӡ� ~)�myo�9+P�~�!��Z�̴�n�X?~Nz�O��_�֥�S��ʡ�����+��7�|�ꑙ�rƌ�]�ٮ��}���߃�{qN��Jr��T�^Z�Bw^T�N/A}�L��:/��X{��0�q�;�����������
2���:����T�ɬ�J�\z�0E����w��\]�a1�E,�C�62���Svk����d/�7i!��B���ʎ�<k5.}�?t;6��<�m���SL��5 ����;�:�G&��W�G�j�G`#����|��U��{^��TB��0)���&k�����mz$�N�Z�I�0hm�����AE��5�8x{�@�֝},Ϡ�R@�Kr����^���������I��sJ,��NayAԝ��Bqz2	?�� ɯ�B���e�t�ڿm�34Oɢ�P)q�Ęg]�0����u�ߧF��9��Wn�i��?��и���>֗�\���v�ױ1�������[��wd��ԟ�_~���s^"�ܷ�:an����{߸��K%:4̜kxo>�f�*S��t�g���1�(��b>�鿚*C�0sٺ.dG�丠]H�С{{�QXh��v����i�y���*�6����MC~��=�/B����.3�o8����&�c��2L�ֿ�Dd�6�`�4!+���jk� ������mqp�XG���*��}i�d�Bɑ���ς�����_c�h���dwW�-���Ps����e�|���'���P'��jV�>�'�6�C9}[��4$�1�9p,Aԫ��{7"�-�]4�I�Ƽ�B-��@��+8-2�����l�|Rd*�H��֥�L@u�á�#3�Mgݖ���_��T�JĦ���¢:��l��4�i]6~Ѻ:�����˟k޽�ʣ�8K�%~�}��;��Ct�|����#�VY�VxT��Uf�e-3ֿ`{)��2�#n�؆X�WV��5�>|�\�-=�0bՀ�ҞAQ�A�9�7ϧ�(�2���d�I���J���L��ǈ�<���l+?�QQ5���5JV���RS�aJ��{���VZ���[};ˠ-�b:c镊&���z,�0���\��ǣ�є�sYh��֛�����_����c䨬������R�>���۝벗�?h3�F���[+SŞ����rh���	��a�)H���I)x/��L���2�"?�A-6n��m��A���T	�2����Q�	��vދ�@�}���l�B�+7�w::+g[�չ��{k��i ��+�DC}�f��V�-��۫Ӏ1�|*?*!��sa��FP���3��U&�����`��&%e�mGr��[�m[+w���2����!��G�>k�t!$١H�����J��k�q��>,�W{ONk<<:zlD2�_�ONz<���Q�Eg�l�JsO�[MÎL%b��	�߰����b}WE�6�y��_ف#�� c�k7�qm�=���I�\�tG�[�����\l�����ȱ���f�V�S����!gக�Q[���)uЪ.��2f��9_�#i�^ tJ:LQ�_�z~�z�'-�=���vQ�a�xRXR^���	����shR�)�'kJ�Zs��l[�[�V]�B�1益q��f��Y���c'�.B�qK�q�����@�~��!��DEE��}^}
R>3�yCX��j �V$�;62|[�}�1^�N/C�dVOZn�;Z���lT�I�R�~�?௩YA=� ֨;b�T�΋:��V;$��a���x�j�c���k���p ��<A^�S0zCO���ο h�:�@�Fq懚�H򞪗7Q(���S�������T^j�>����D;�̊���b��0��Jl�������]><���ׯuUK�D��Aĝxhp��ߪ! tԉ}�+߻Rj��j0&�Zl��;]!��5���m��^�L?2���}rv�:U��3�Ώ?�t9�!2�Z��(\����c�Y7�uJ|�)�$cha��)n[�I@}�"9x�����4�}J���Ҳw� i�DD|�󞙆a�'%!q�A��Q/�G�1�sko�.�ϋ�v�C_��O��]H�tSUQ���nd�Sz/gm�Ĵ^�sl5������.'��塢$,�N�K���\rg�3��^ȝS���Qm�&[�$s7����7��p�8����JKqj�����I��b��󬵋T�l׋�n��7�^��%Ϭ7%��ht�Rʕg{{�|��|bb���s&*>�.N�b}���#Y81F�D��3<�)+�K4k\�ݴd��cK��-��ap��@%���Gy�� ������m@5����Z����-Ό�"��~�Y��c7D���ZG�x�W;c���ks%�ԖhE������D��"oCV���#y�V���C�B����a@��C(�CD$1\�c'Aȶ%7yu�'Χx$n�6��f��OF757˫��
�6�U��w���n�cm�u�v����-�J>�ɶ��[���蟲���s���C��H{��;���)�K�7��f�ұ��@-\j���a������D���p�����[����
*��ʸ��@�+rr}��t�b��z���Z�X��Y:��>�q�k���_����ҫ�fC!�'�ɯ��LfZ#��1q("Ex��� �tw~�Ŕtc` �4�T���o:cd=�9�Ix-������7�Lx���o众"�Lx��gT.wVt���i�o4�^f�����2�fY>�5Qri����O)3"aI�����!2�K��4��O�!9',�`�ۘ�B;>~(����W�Z��X��g�:����N�+=��	_('����u�_�r�����*�q0��j�N�l���L[M¸�Xdx!�W��i��X����1�xZD�T�}ڔt�����Z�a��['�#"zt9a�1����wO����_��������<`hQ��*q!�	�P�uz���A�	���(��W2��˱�DJ�9Jbz�6A6�.��7A�|i/�SK��$�/VV!M=��ڦ8��[��聳8��/�s�4nwW��f��A�X�l�GVm���<G�UC�`��"�1J䎜`��^������E������s�%r��݃�c������}*A����y��ᱵW�匛���8�=���M��[4�bB��O�f�v�ȸ��X����=LB���;�"E�<���M��Q��2��3K��,"Da���ת�p��.�����1�f}���TC�>:�uu9��s����2}������սo�0�#BEO�A��_/�
e๸�ʗ��S�a�ɜ�O8�VGA������X~������_��e��yWKF���a^�j��i����>��d�݇2An�&��6&/U�����7b��$�x�(�B]v։�tE&�z܄a��є%�fk��8P����M�{{/�S��z2%����u�mݙZ��9>��������!^�/�tGh$�;���W(nK:����4��cf���Ϩhu�����Zs�w߼����We&�$u9�{�~?��?�y�;(RvͻQ&���Ġ*��B2���T� ׼~R����CjF��DRa�1�����<� �C����.�v>�eOF�l��9rˤZ����1�eETux;������m}��[�y"��e,�j\4��HR�Ϙ3UV˕������7����FF*��?��,Ty��eX�6�ݹ���r�x�-^h���EK]��	{g�4�Xa��@
��`����g9��HG��\�рئ����w��CO �c����&��?���جY�t=�W&�m�����)Lm��\���2��^��Cȓ��w���BB �#C�m_�NLA|Iu�YmXK��z��e��o�[E���$%��0J#[�=�ga���z]_�:�N��S�K!�B��a3���MI(����o���}�����3�G�d%2�S���.9�/�T~Y$�$a�3x��HVL���Ցjn|���������ֽC3��҇�t9�LTP�4���J9'�:\��] ^��p�U�\�h)u��,�����5�"Gw��Y�cs��,y�W���SD�(�BW'��|�v�uǋ/&�}W &}_3=I��3ܖ���؃6�fe���V�Lk��_�@�a��Y�Ư致ȉ��������kyE���^�S�3a��>lz|�5Ж���]�������^̓fc����Ek�'��� ��G["��@�C�|����_kr�&aP��Eo�ŷc�q�[��;i���>46�H���RsW�<aէ\H��4��R���5��ūF����˹����끶���N20�>���s�����KA
�0���7�f_�`�	�z�Y����O
�?w�6 ��q� �~��}F��� 7�k�����Ŕ���Zc�~Ԝ�f[_z��tjH@8�]uo����V5����m���́~��y�&������w7TbOL�*y]x�=�'��SVl�U���ܸG��Q�I�,Y!]F�e\T��m8	���S呈/��^9�9[�1'��)A�Q�qDs���~p{���b�, ���RiȠ���؈:�=�3'��U���'�y���'|nO��r��7��,	yZk����ڟ���1�$;P��������~������"��PB��c^R)�إ�J0G��̰�5��x~�=�Z��+P���?�t���������K1%��Y���f[ķ�Kp{\����o�����7�4��y�H��^[h��\[uINX�w'���kC�ܩ�8Y����;�f>\V�wg_�F���)-�J�+Æ����iR�Kݟrn�~u�2/�������rg�L�k2ѳ�v��4�]�����������v7i�f���=�+Q�F�ë`�38�N�͠�r�e_��nM��\\\��7b�U� v�w�8�<5��zx�{wC	���2'�-�Q����o|M�r�s:"{�����M�v~CCCe�y�s�L� 1?��2l|����i���L���������A��2�����2��4�k��/����a,�F�����̣/���)c���]��^>M�t��Mܶ8�*���v�&=#���_w� 8bg5C&dR��������z8<�k��� �(n�hwo/gL�����8�o ��z�#����b[YY�06�͵�ѻ.�cS��=rZ�SY?��^	��&k4�\�斾��������H[��YC�@8j��=������:
f��s���U$/T@���lU%$L��Ю�&�%w�S	���a}�~BO�S�Тk��b�5gв~n`�Jab:���V��lsNG���ѯ��y<i
G��t��@�I#�4JxTh��+v�gg�+�KI�(���QS�^ۃZ����@!I�b�h������f}��3�1#iD�����\�:��8\�pBZ:�,V�d�v�����ڑ�}����2���Җ���t�O7��w��鶻6L�8�A�A���;�],`�~ΐJ��Pt����������i����^v �)f�y��(� �;��F�UL�ٷ^3����}o���	�(V��4wtT6�8aV�.��,���v��������Z��\Z�{e'���L*p�K��T4��(��b�������ƖS�� ��B���W��A�YBrZ~��Ď<{���)Vl�{�~���a���D�"�+m�s��n�@;��%��%?}��x�čLZ���I����&!^�L����O�XΧ���D������M#�/�
�IC��3~$�P��|��� K"��m�3ڶe6�8��[FȒ.�Mn�~�vsw���;�s9��O#�U0A.�c\Rw�/�!i�#�7�=���i�pp���Z@Kd ��4��4��gzi!�bg��u�9୞>�f*�˳q���U����mq@��q��	��?�fe)8KxKgQ�3k���鼃#})��	��-`���m]v�̤�d&}h^wy烑�ߔ�Y�Pa&I�23�-����wjl�)u��L����D������c�f��m�О��,�=M��47}!������=�=/'�������M�ƅ�Z��D+}�r�e�gq��
G�٨5��:��a-ψ>-nd(R$�|xI����=�Y?k�1�\27[��8P��_�����h�}�(;nB*� !���N�lh[c��O�U�q�I\-N^�V m#�DU�>�UD8۟�q��0�w�8���2J�����
�$�/���<�7s�6����N
�jJ�WNl-ez*.��y?l=��F�i�=�7Gtv���<�tWc�ت��--z���,yF)C�2�Ӂ����͊�@�$1?����A-`x!oѲ����8	��/jf�)�w�g���p!֞����ڡ>d��� 	*=
�}�!w��0x���:�_����+G��lEx��~M����egaꐉ��p<h������+�	ny%�n�0��w����l��Չ�[��q�
%ыϓ��+��J+I7�E�"�e9n��h*�o���>���e��f�����3��*F&��7�X��0mƴ"C%OD�"&	�'(Q�`�,�mN�ۭE�ׂ��ܹT� k=��ç��&^�`c�ڋ�Z�r�K�H�h��Z�1�RY���eR�!�3��k��v��j1˅�R����%/��)����6��Y�b�=��K���W�y��؜���$@n�;��iŇß��KoL�_��ˊ�?����7ܚ)HIKS�Ho>�BWS�^����쿇/N�'�<:}i�5W�~w�������]E �x��$+o⺝�F�Qpr͙��(�=��T��&�`������P#���uĞ=��d�1�����No������v�[��ZUX�~h�������k�� Ik����f��<�Т��9�k�����Z���t-	�dgA*��㬮4[z�� Ő�f.��k'g<���,�V}:$��B:yp&oǧ�V������VZ�h�8y=~��/qSաW����k��H-97��2vSʪ����{�v����CCٕ&	����SN ����k�,���l��WF?����1�N��Y���e��a�b"�)��O�Ɨo���������)���;	LH�1�+��A������BЎ}��b'�v]�>B�u�),�xI���l����㻻�oT�W'��э��yx�����f�J�h/}*�ׁ�����ɥ=�P�%�4��@LH��	��F�S2k�-o#1a�@1md���� q��OY�vF�_B
'@:�W"7�+���a����W��]O�ܞYܿ����z�ក�'>��;���!#�d�ћ(v`��X����%��!�Q-=������S�B7F���b_P	�`������&�x)T�����Q�QU�6��/�7�\^֎#��Z���h�\�=�1'q����.�<}A��s���;{D@U��:��əv��o����a<��i���S1]˯��H �X����+���KƊ�qc�I�Je�u��Z37=#�x���k�P����R�z�Ȥ%�Q�f����yᡛR���!G#��T4w��tD�?�������.o����/Þ�}�x�ě�&��{]E�a�Xt[fr:�Dq��eUf���.�����C"r݃��V���u�Qn��鴄�.����.�AZ���q�9� �i z�Oj����$�.YI'e�ǋ��ӝ_-�ɗ��}��	�l�Pd�}"/8�u|a�в�dZ���r<q'���n-S�z�'�����e۝k�~�ʹ][�������뉬�a;/��ƍΠ�PI;w��>ǭ��12c�q��J�^9,I��y�c;hׁF��OLW�����L�\���)sa��-��E
���]��7@�JY�ښ۰� <�1y�c�K�0�H <��h���t�7B��7U��n�Ϩ�@����i��0��g��N�>F��~�8��O=����I΁XnY ��.��\>κ�\�M�I�.��CM�e$8���g�=�"�7[bo�U���� �\�@k9��%�Ñ+�[6�&�{3Ҝ)�@�֎���`�����;}30���{x�sܨ��ҠQt�jta��&����cO:±'3���%���@O�s􆧐�p0��Oj���yX��F>��&c��'������E�0n!p,��+�qx����ȫ�D��\׭q����ߒ��-���ȱ�tp3:Q��o�!N���Z�Q�o�Z��Zp.Կ&�S�J��*�A����e��b����H^�r��Q3�8.S��A	Kb��?��y<��{�\W�D򒢓�h���g�' {�v+���=�ITa�����Q��&::А�뜂�2����O�+���z�Y'��Ǎ��G%�P̿�&�����2�u>�����{_��fs�'�ڮ�^�KT���?�ta��ׄBe��MD��%sJ�2���߶�ʖ��7�	ATJqqBC}�b�
{�BI_k��،�W�%�F���D���IO4na��7��9�Ҟ5�t�Q+.����"�W	!}#�gz0]A�X~䧉�`2���� �泀b�]E��qg�E�;��3K����P�l�%1G�n|u��)Y�>���B�-����{P�8��������Z{�n�VV��.�dJ1T�'�8(=�i�|Ϸ�cN48��CG�H�!*
�z,�u��L�u=!�����*�b��'��ɑ�]�.�&����*3�(�i�A%s{t�����uW�P�;�_��$
�HeM|��J2�TQ �?���ԕ�}��!��?�~�6�Ϸ5��x"���ɬ��!�if.Ш���I�����
?	˹�u�����`��t�Χ�Oy�c$uI�F76�@�oM����%Z���}��U�$44xҚ�(�Ç���zߝ��÷��`��LY^��ȳW��=|K���V�L�jFvw)������?.������+�������s�g��Xh��4�7�ōr9�� q���p�d�* Vh��kZ������Ϧ�y�P��76�ttj^�� U�6��a4�x~h��A�3)'��X�<	/c3�q���3�t둇�u��Mb�5\����X�6?�$*($47�+�9k����=w��6v��գduBB*����s_����7�G\�ZO�����z^7;�(�um]��7N�ַȔ�j�I�~w��!���~k<\��LR�j��F�O������'X�[`<U�1�8<G2�Ϩ�F���J	��
�]�5*	p�WKOW�R)���gԉu���6�hi��T�˕�����Ɇ�@oP@S���8�f&��8�Y
n�d������
}p�b����|̪~\��^0���$Y���cϕ0�����c�#M�Ӥ�E����`��Czq��������žag�����	|�g��s0�^�v�l�7����p$^���
�,9#<nJ��}i�a"}���0��ރOpٖ�L:�2T���	����h3��U��$kG\B�a \�{ X%�G6��mz�s�(@p<�|�X�; #�_z�����������i���H��ԭ-��<M��0.7�����FwLt���tt�e���JwkJ���m8���<�e��iK�����P����r=RB܎=�Ƃ�-C�ĻR
�C##,SNm}�'�[H�����/���%�xӸ�3e
-R�\V�:.�D�3*\U��B7aG�I/��\�h�8�0گ ^��aN�v�4(��qA\T�S�=�V�i�( P\��:�{_m>J����_��������Q��o皽n�y����o/�a�..S��KA
ϗ�I-0r�h �����~=Ka߿ĜB ��#�~�ׇ�.x�-�N�� �^�9�Ns�+&9��>�)/ %����.US���Z�xFt'Z{�/�Ʒ�)Q~\��z��XX{pl[?c���\Xw��dw$�~5�Tщ$�:F�w׻-����`��	À����qF~/���W).�P�c{������H	7���M,���!����f��]���P*�+/�����\8@/��m||�RR�c��vw��j0�((��<:��^ȴ�l���k����\Au�Ѣ�B�l~��A�e��]�ǐ(�ӏ\t�v��	�x���6k��$g(�VNZ��Q�v�X��s���<���1GϪ q\V\@�,�>���Q <�[!�����Jhn�`�B.z��h�D�d����: iI���~�/͍߅�X�v���6��;	t���M>)�տ�8�Q�)fG�8�ȝ���	7L��L����Y֥:L�$�f�jTd��ΪC�@2ɘr^A5>J	��5�&��|x�c�K=x�%h�ˎ��kGK����>��m����V�+}E'��[�{��.^�� �Z�?���)�����s�|pĹ�/�:�om������l|�BăD��t�N�勍�(�g�'����J2��0�F}�2��+�[��T�BȪ.�s�����0e���� y��~�4��%��i{/[EP��� %���6mq�.iDmGF>��0%^�2,gn�#������8E�`��ꚃ���Йw�4�̒m���T4�ޕ��++�BY������9����	�`�p�<�{���N�́�/��D��^�_ܑ7�s����Cʷ�ť�;�p]#I
��9��a����Ŀ��l�#D�Q�9�4K����&�Ƕ�r<�r�S��?!��{�{+?g�v���Q���E�~��Y�����R�"S@��('I�f��ﭽt3Y	�p1�C8dV���ez�6��o�E֎�<���0%��-z�*�[�N�]�d��^�.��f����u� ���r�����U�ڧ=�3!����zb��Ei:������U�L/,tV�z#� M��LA�-�]D/|Z��A���>�-�#3a���kw�CL�f[s5X��o��y�*K� }�͍��a�]'�����%�/޼�"CS�Y\��h���+���Γ�o�\]��\��wS5x@ 0圯�Lu�&�=�}+M��{p�X�%�p}C�vF�e�_Z�柗5Lӂ�7���U?Bڰ��� ���mIr��~J�������m(-��
��L�PZx)#�k�Ee�������nc�e޴��o|U Ot�/���'��N&lqNLL�Q����:uW��hc4��������i$�~�=\��v]~;��?tʃ'
�VA�@�����V�܆�l*��V:m�����$�]\����6�ŋW���>IR2�n�!]�^ihJZZ�Ėzhy��BJJ���)g�_~t�@O�Aoqz5�79H�H�n\@c��Ln;��[h�Q��B��N���6���A|����-�FX���d�g�^�����ǹ���@%F�B�O������i��N����;����WCC��	��f��2M<�|M:��)*gOo/�5��������^��{zF<��im�V+T\�	2��:�/�<��2����x���LgOV��aj��i���j��1/~�[xw���M��#�yFF*��}���i���y����X���~P硇� ϣΗ_����nȗ���Q9ݐ�����P*C���=#Ԝᖺ�b(��:� ti�rMٮ�y!�����w�ru�GA�%��݄�c �F��ͻ�º��� 
k��X~QE�}�˰'�I�\��¡�i*�J
�U5c?á�5*?�� T=KN�J����}N1O����ϟ�?,�ߟ����
^__�F����*-]-���5�M���z��jЈy��DsU�����+�������"L����6C;IC����m����5�PpGDX���(I�ۺ��%H6�3�,933��by�|������#t}�H�%�*K�y���`F�D� h�hTH�:�G�K4��ꭄi���5�4?�* �T�Lh^��0��[�ҥR��t��S�?6>zB �9Q�T?e��>@�GXn߬���G���ԫ�LpK䪘r
ss�BkcLz�^��c�E�W�U�W}��*�r��J�W*O���V�}_sxU���󦠚����	Um��@lg�)Q�i\֍�g�T�w�ݍ�/
�ۚ��G�ݬ��bG����j�A�h�W����#����~[n����d��#gf�S]�QrI f��M�ɧc�Q(��13�4���s&�M��0�پ������y��C�C������S�m��@(ɼm��Ӊ�rR������E�����h}�+�z�T��m����[H{��;���P������N?��_-�l�4!�e��t��>��q��U��ZGM���(qQ�V�H�`�_#)��!.M������x�[=|G��5�����uP? p���m�����v*}��a�L��"��w�>�� �C}�ɿ������DaKۥ�=r��t�W0���-{q��=^������kwᣟ�����������L��4�Ob/�6i����ml�Y|[}}aC(-A�Q�>3�9�&��OK��9�Xl^DNK�5�E����1;��k]&U堏_�ؽLt9�7�~��/uMp ��[�C%ȭd��]]���6Q9�~�����:'ЯAиD9��9S���� r�+yg��K�"����R��` ٛ�Y��`Λ�����o^�������3�s����V�>����|&�-�b[J��w�3�˗4���oj<�eDD���V��
���L0�T��'>=?�(%�YU55�2��YYY���$�9��b�rt��5�뺫ղ�(��C�ss��*ɼ�3��h�lC���[3N�e��m1Z�XR�����,m�Ķ�6�A��������8��˛�ƥ�>��$�`l�BB�8�⍥5�I��G9�Q6m�;]��Ћ'h��B���0�������ojg��K���y��n�0]V #�x�����<�j��l��A �=y�3�ѭ�Շ���ɷv�ߖ��hs���٤�����㪟�jl`���u���*;�=z�@���C���:g���FJ`����ŵ���8J����i1ql��-�פ���ؽP�?��m|��##�wԑ�	���������8^݊N�E�94���e1�58�7�G���o�y7j>IL��b��8���x'��g��!8Kz�[�����x4[�e|J� � 
fDO�D1Zp���^ ^��<���Я�?H�bv�1~_o���s�l�XiN�C8\h �\��!�k��hz�TL��v�㚆��X���1�ml�||��C��K+E�zi�*�	���t�>|�M�Љ�ؒ��b#�b[��qȸ�ԃ	R��#Y;?]�Ϭ���9���[�|S8�&_W>��S��o�wOހ��L�����ו��i뮦�l����DE�3��_V>K��Ƈ��e����%({su������t����(�r�2�����o�Zl��cFk��e�Fe2�Q����ݡ/���ޙ��6|�yi_��X�@J��6np� �1�!��0���w��J'�7?����FU�<�������;�����7oG�f&��'Q�n,�����܉��-�3�l#�,vv����32l���h�b�p��ٓʆZ54��e;��N�c���* t���YX��SD0@2w�U��"� �G�h�1 ]������\¸[��w����1�,���/�)�%�d��c��z
Y�J��͇�yK0���2v뭦h��
Z��la�%ȧ2����d�����@�lQ�ޕ}�Ճ��c�6�o?��\��]p$���\;�0��sj%f��gQ�䵵�]NM�ii+f���92��pdOw�Og&E��"BB±%n�.��Υ��Ƶ��~22z3�0���RԠk�@tSX�־�>1'E���/4j�e�I��D�)��w� �ƛ􍩫O�"_��1�ی�V"±��!ׯ�����z��£b|!�&�[�⯰P�o�'�v	�7Ϟ|o�̩��<?��v8����o�WA��c����&���a^���g��̦@��*�`�=R�~�Ƞ"��nC�������*|F^Z��D�B%�ϧ3�6��a��Sų�aq��PPRb�hw��]�������q/�Ȅ4���ޢ{�㰼*J ��77�/��+K��EKH�`��ԣ���>���_͇,����⢐\�$���̬:^P�|=�r�
���\�w:(<]Ōn����@���y��b7�;����L��2��t���䲶���-	��:���У���2������O�J^����ؘ��*�̳ܥ'�`=�r֓�M{U�ӟ$͐8�s�4�&��}��f�<�����	~���S�nA����qK, �g������ $�"�b.���3r�6��5�"Sh)�Q���x���&/�a�!͐�o�R�Mr����K��Z� 픬N���c���K�Ӆ�q���xC���g<"����̥�ޒ�[��S�9�s��,S�D�1>�2	}o¡� .�%G��{~9�r�n�3�hl���U�D�V�������E�$�-QC��H i�
?�4��4�Ӡ+K]�(ח�ڪ�'�崯Y�ig+��h��`���^�E�=sbUus�ȣ�:i�a�0�xv�ܞ$g�ɵ���fa��";{�:.Z{��9��4�Rє��Qe���%$�&\�;���~��^�s�o���8��&������Y���lL9�/y2�����!��
o�
n�����[��/�p�|���V��r}�ґ�Hʾ��hn�u���Wc׾��1�%}+9Z:r����⚠f����tvP�2yc� �k�'i��;f\�P�MZ�h��}��n�({o�A����vTK|�7]v���u�uB��u`���k}*ьP06AHLo`i� m�m�7��C�� ��3�2��Նy�^CfT�z���ң���wtFn��[��&���D,��4�'atfI1��u�QQ?a�_Z�I]$�n�%%$DBBZr		X�DJ@�KZbAJ�;�[Z���<�{�(�ߙ����\3�]W�E_�f��|���ȶD�\ ����n��]�n��Q�v��I���R���!��d������^8��cWQ��ǚ�2sxA����3�E�v��H�m�9+h
E�1i8m"�9v��		؞�Ab��;X��ڕ�CH���3�y�C� ӪB�c|<O����1���ߚ�c̴p�w�}Yo�JC�`j˙�c����1����y��L&�QaJϚ�p/��1���e�z���=}0��3'v�e��m/����R��ba��%��]���&��A��G%7��BE)\ ���ippmK��ԩW��#���ݨ�/w�w%(��}��$&z�Cu�d�{c�!E(�OZ�QK�(!&��a���c�<�oW9�$RTUk_6��̆�kTr�k)K^E+�?�9)����DT?E�*���vo|����R\�E�h̶wm�OZ� �D�Ҙ�;�r�D�!zC�	N��&�mrqޤq����[IK���Ӆv�|�&��As���p�
j�`��9��Հ�7��t�h��[���G�\R�9KMrJ?0찭(�0?���.��;�M ����;<��r&<��)����x�s��G�cy����{��N"�W�=�>CNL$O2c\"���Ӭw-�I:M�W�~�������H7��c���y=1�P���ƾ�g_��gT���d�>O�W�I�߱�O	X�9�� f���>��� �Uv�Pٚq���xWUc#��*���oݞ/_�v��������֯��J@�5�s���<��7o�r��EAFI AAHXX��tK��/�{��c�����'����N�>g{I��1e-�9��JKD]*C��<ٷw�Ҩ]?�|v�]&4��/�q)��%��F���D�Ndg_��Q�B(�͸v湔c��l�V �.,0�n�%�p��ؤO>SP�ǲ2�.��!��+e�� i(5777���ulfi9�~~P�}'����2L���M${�g����(��T.w�����
A�
�Y�v�_�N9���ۀ��۪�~m�"���Q�YO�S��8���k�q8��m<�zG�D�t{�2J&4��D����{���N�6�@ ds�}�B�ψ�♒��1!E{�>���P& ��)�2����Q���Ȯ�%+���4��r�6-�%�1��y?ŉ�2_�޲����h]�)/�X����8�n��(�7�	�wj��5�YJgfga���2�^߳�x@���R	�=��P^U�&�P��H	.]T��k�f����Ƨ`���'Kt�1�`�_�r�m^2d��ߋjW���Pr��w���o��nR�J��.�Z�0���l�F'�;i��Q�K�(�Z*��D���|,$j9􀗊�a�:WF��H�>&��QfJ�#I��H��F��咲�LN�	�4uC��K���%�3y���=c/���pv�5��Jv����@*0�����+�^�l����r�6�N�I���")Ca��/�&��l�p�;Gi�P�W�ء��ѧWZE��5�-l����V�?	�d�7:*�:��n�Z,}L'
`��~AшuRr�YQ�yΕ�$�4����aGk�x�Yb�<�6FsQ���L$��2US0��a���3�Ӕ]��;�|J���ҵ�11�6��ٞ�uU�:/?/���hD#t!��P鿻�[[v�Ҡ'z,��o��t�$V�u��j<�i5�hm�Í��}�ȧ��1�a�]�����C�E��S�����wp��ơ��.H��[yK�Bm_��@mc���mFA�G�ԣ���S��4.X��9��;\��/(e���k�|�~����$����m?�&������K++˷p߮�G����	X���߁����K'����^�Z�'���������%����&��h-�.��~��3�fŶ������E	�y��Ml�`YDI��0�"�I���=�c4��C ��Y��YrE�h�F����w���衪�ji�K
=HՈ���U���.Ԅ��E���Ⱥ-� �e���R�/[		:�~��b�A�h�}��y�Qe���e�Q�`�ޠA	jgJA� �6�3kM����p­��4E'R�&���������bP-OtD��z�̩q�V�\��17Q>�ΐ�_֔�]m�<򩴁�e����+�P��'>������A�U-c�goZ� L������ww}p�d`!�[f,}��G�"Zj���da=�e�K.�/VɅ
]��o545K��ZF��"�e��R��Jn��&|Z�$QkV2)�*�q
D m����DA�".����HH�Q_��5~���QC�u1�q�Ä�9�禦�Kt���U�P����v�gtyyZ�T�ޟ��百~�j�Pw�Au�9����R�`b�������S��L.��B4q[%!����[C�ެ�DV������a�� ������V��a�gZ�ӛ��wH�y{�����Eӷ���q�'Hě��C�-_�k���1z�T�3W
��!XwzS�eC��'Wwp�A�B���Ώ�ص,�媃��zlO>2I����U��W����H"��@Y�Pv�G.xsx� �&�e��qe����C��V��b��4�v2U��$6��fX�ǲ���G�j��S�}2FrF�������|�&��f�4�����]��$�{n���B$��b()�xDד�G�_&�5`�x�� MD0?�D�Pc]r������-�����±7�<���[Z3� �u����{=�����1�S3�,�E�N�"N"u��h�q�Jѡ�\8:x/�F�1>N~�2�T��Di��������d�O(8𿎅���!Q2����{;mÀ��'���-a��ꊞ̒��48�yg1�ț�B�G�}(Ѯ bMJ����Ev�Y�ŢuA$#��/����]����&eT�1x�ٷ�C��u���ͩ~2��sϹB<�윃�߄��������"�i����~�<<mX5�p���p1�N������St�!/��J�ҡ�y�B�ĵN������q��ׯ��ЛƀY(�gs%9茹���}���(�rI	[B�E��||��hA,V;��x����Ϧ�zy��I���5� �-��\Ӷ�A�_!��"d����<�HT+��I?%$�@����L7�@9�v�H-�8F�7+�0�
HJ�q"�Ǣ#r#���[�K�r��wα��[u���xR~��Y|�
��/��4^9;+�~�f+�U���ϒ���MX>�5������D��)�B�whg־gӿ��j����!�Z4���PoD  �.�%�.������㵷�P��9燤���倮��T����8������+�� �.���nynn����6x��*Lr��4���q�C��=��Ȕ�G�/$�+����pp��Eޣ�a�N�ϩ��ٸ*����~̐��"��=�it-�� [b�n�ǙP��es�3��A�[1���y�� ��n*�|I���\zx�=�7��sŊȧ�q�k�M/G�r�1AP��	p�؀��#�f��lC�|��&�g��cJ��kAI�Rܜam�k���t��+��췹��mx���y���H�����Ŭ	4����I+���ti����uw�^AUg�f�Ɔ�������*%���z���)&�<$y��;��a5Ů�i"`��6�p�۷�9&�߼y,8�}x���R����`�V�)@�{���q=�A�9����1~�Cf��3Kp?�lk�t���5���ݴt���ca��g�N��EK�D{�gr�4�Pw�A�L�)�M��D����7��5,>*d��9C$��� �\b�i9�P4��)�!???zgǝ��{Sn.9��#�����dƥvV����m��шU��	����v"���񼘥���T�V ��e�l>:q�X����������8;NU=�v����_z@8��H��B�
u<3C�!���)Sh��w���~�
�	����P5z�?�lY��~{�4�>�a'K��� e �ɩ)&g�啟Ɏ�s/�p�`1
�˷�9+H8:�T�����4���(̴�2�\��bm i]�{$a�GW��}p
��q����3D]�C�o�@�G�����H,�ǯ��sQ
kݱ�N������[�5��"�ìպE��[dq'|�A� ���N��-h�ꄾS�&��$;f{�O�����x��K<��:�~��	��"ɉ}_z�$�� d�@��L�R�����������@Xp�P�wꤪ"_� ��ީ��ʭ�ܡ���R����%)��u���� ��*�#w0��
m`P2 I�5�.d+./�sQ[�k(Zt�b'�m���f >&3�j��x���(��x�j��U��ü����0�qt��$A�ĹR�G �${�4WR}�Έ�gC-T?^����˺�p�|B;٨�vV��Le���>�z����Q�)��&v�����(�'�q�+�ٶ��߻ s��\)>	*�9���Ҿy
�#qO5�fgu�N/�@�2����h�JH��ZT2^!{fgi{�}p���!�pi���A� t���'��	��ǣ/�gR�@,���4Qמ��,7(����`	dc��W��x�,������6e��e$N/>��A�Y��g�B}���]N��
��;Ƹ�^�oǗ�?�[���\%Ʋ�O��y'��a*Ùm�FMNE�<������C��U�&�rƿ��T�(2PY�
�%�~��'�Y�5M={J'����'tx�Y�t~(���1�K��a���!M(�����ɿm�슺:�A�����yh	�h�J�}��E�@g�wS"��q2��1�~�������w�Vm��5:�<��wOMLA��:����}}�f����ڏ�1���QHzz_�`���)^%��-�}-�Gm{OcUa�<:�m~���ڿ-�_l���c�J�L�]�]���0��a�����͹��J�����_��y�?j�F3Kc���ҝ����=̿~���� �L���������ӽ���k��;���I0�f)9���=�P�B42�صG����u¡K�ّe%�,Mu}�u�\y�uC5 �����~D�mM�:`>�/��C2dga%'�h��C�h�T����H�5QL��Ԋ�3�,fh&�kFhH�Q�����|�`�JՔ"	aYB�!���e�NGO�(3�3��H��X���Ã����,�I/u(�H↕���L��;��Z<<W-@�u�o� #j>���q:َ�ۋ�s6�����ϙ�����{6u)�J�b��S/�<i�{"ԗ�2ד�gO�qN!3F�"�gͽ���H�A?�G���z������n�����X���7�f��;CI`��R$!&�}�#��5���,���|����ÿ}A��k��BܠB_K�]J�>���|�Ƅ��+�0����Ƣtܥc/��N���EO�HJJ"7p��=�&T7�0�� `V �Y���ȍ<�o��x������:ߠӜ����F�T�F֐u��Q�г���^
���B��+ߕ��~����6�����%��b�D�O��?<�:n��b_%�����,�da��4����A�2�?�D;�!�"�zN��l���w���e`����!��sX�ݺET�75eLYO]���j�ϩ��C�iF�r�y��Ą�ë*�� rRO�%�q��0���S�D�^^�G/�n�_�\"'�:��Ѻ�Ǒ�W�j��a�Z��c�_��r��Tw�74��چ���e 暰����E��0Gs󜃩���ة�Ci\��ӑ(�D)�q�Ũw�@�����=�;}�vƺ�/�#��LY=G�D;�G^w�տ��zT�2�E��^�Y=@�RlA�X�9m��Bv��mܴ6��^����G�΀�����zc;�_9�}�w�� R��Lsy3?�o���z���2��"����G���{�7�U��G��e�����GJ���7��˦�W�/O~��T<�������53�.�3�ݽ�?7�1�V;i`d�owo|2L�|�&ܮ�gX�5��aYM���]7������*-7� |���Mئ6�κ���Y�� ���������u;�a��n<�鹈0$����$��(#���yP,*&�ے�O$� �OD\\{Tm�VГ��!2&�n��f�)Υ8{e0�G���1��9���U�`]/���*4�Di��B��(=v_����DuX25�-�}~?�w.�*_�t�|���ҿ�^�dT�@[�4�â{#��bLp�0�#ͅ:F�6�2��v�,�@��t�w	�k�HS��_��*���v3�%���r���	fk{;!11���J�j2�e��a-)��<uH�����u�}��ʦY�L��Q>8rG�9�����go5ED��쐅"���So[W�܅$nm.��ٸ����4��w!3�Au�����.i����,:h�khK��z�� ��d��g�Tl���c�^����D������Z�.�A�7*���٩|aC����,3'�j	.��� ��O�SD��0�=E�^GS��=�G���eф�oOt��\��1�>����Ժ���6>>�/�)�x��o�S"���D�����q���G��_�����&&�n�F��NN���T����P�a���
���˓���j�C���J5�i]^F*i
�<֚�H��z+���<~t�\,d	~85�rU�[E�c�I#:�a\ҕ�^���w�S��"��n2���\�H_K.x����Ѯ�꘩uܿ�9x�9ã�1+��j��S|6o�ϲ�]N,��#�6������j5V�hooOQ����sk�TPޟ�rs�'��s���� Ǩ��&T[~t��[�w��[��;��N��4I&1���D�����TUUU�r�T���WL&���h�p2���^)�T����{~e���cCm���^��p�X��ؽc���Be}CP��Av,"U�Ґp�Q��'������j���6��C�Vv��d��f�Ys;�"���q��۹o|�ds�<�Tߥ���M�����6����\�y�9#6��u3�J_�i4�m՜٩�C�t�	\^C(�`z�l"RRq�D����;
���HC���%M�36rr�E%��� @����vya#�PZVF���3;��9�s��LU Cze����X�-l�v:������4�L�j��շj#�N�L�����k��2��X;Kxs0�m�]XmU�8������0�'� p����ё��津�/�f���yI{�qs�~�"���7"�ƾ�fe�t���w���s�@��8�8D�E����ͮ���!�-��$M=NHDt���٨fEM�����Tt��}��	�>'�XQ��N���2��@lni�`��M}p}�rE�g���h7;?��jJg�,2*Jy�1��T�z	�^ѝ� �Xni&S&h�*��^J��O ���J�&����\���r���#7��|Ȍ��w�����`��W�j������4ў���U.?��qV���f���r�O�3��^��g�F�����-�yo��E�j�2�|���Y�����뫢-�O�1G��0��xJ�4�]C�9�~^*�55š�q�4����!�8�\u�cz��N�s��@�pZ�� Z[Ǩp�Ow�1e@s�o��k���oY�-���0-7��ָeR䟷�O��lR��}���տ��j�#8a{|痥���z�21��������U	���/��X�D��"��1�� El��-\�B�����p[S1Z����:����M��DDj�%��p��(�*��X�_�tu)ߥ's��I��:���[2Sf\ƒ1@������Y������\�#@M//ԇg�^0f����9dM��xT_|�hf�9'����,�K�p�jX�ƀ�����h�5�tD p��V�ɟ�6ǲK}y�Z��튴P�=�\
�_�|����8N�ԌI�
Z	����}'P���O�p<����RDտ�l�s�_=�9��s�����ί�_��u'Ya��c�I�Kc�@��f�5�@�(��x0��@n(���E٢
�t�ڟ�Ϸ����-�m���PZ|�2f�^A���H�DH�\-�
}�T���o�){�sc�=�(S��mtV�@�YEAA�|�z��S�k�ȶPw!%֥��Ԗ?��^�F�X
�JH���
�!���rk�:�OL|�HR��ud���+2�y���Ge���&'��hL$��E�x��%ڊ�xE_� =�Ϸ��Iwpa��dnnn%��瑸8^b��be�8ii�QMǋ3#��h��xO^mb�����7�P�q"x�{!3���b��ͱc��2<Y���մ���ӻ��Z "����p��_� ž��-���}�֌,*��G��Qn����j#�u��ȕXy4�:�08��9�BL��#q7���)�@mt��zBh���89V��E�P�6�[�4g�kޡ����U�z�v\����%��j�7ul�ʇ�{�:NN�5K���_\x/��o7V�Q��#ub��Qb��e`�X_O*��ulfcs�q�i��ti�2�䕵���������d������3C�Q2yP�O����Ԃ[���s�٩;�*�0�G��������-�;dƜ��bn�d9 v�pg;���n��e�6R7�r}�'M�Z��"�VqIު�A|pi �X�ծ%dsj󌎮��c�TAO0��\��5��w��Y�n�$2���m��>\�-R9��s8U,�3�5x���lh�:�O��HJJ�E��Λ�N�MM5�Z�GA��J��r�m�}�������-,`��ᬭ��F�˝��.�ONO�TA�~��upV����-�y�a����=�+d�P c [�|�a��꺲�6��R�:C�$$����#��C	�� �OH޾v5���Y�Q��sE��ﯭ&�g���V(t������vS�0�(�f$ԌpPr.*+�~Ґ�s�����;9Ik�#E��~��
�S�"]�]ABd+��g�sk��)h����[��)J�aSS/l��5�fjˆ�(�����iiiI�u8_301=�D@c�He�������S�G�X���Y\�~J�Pg/��oQ�,ꖌ���u�R
��N[aDd&t^PAJUX6��(�� ��a-@>p�_{C���$�)�C� �����t��n��&�Ǻ�����	*���b���ʵ,�K�[Ā�lC^���=wuq!7.��Td�*�88�y)��f�����f�-l���!�n!�伀����o/�yh,-'��&dJ�������mG�T11�Q5G::���}�O2��!AXR�#06���	�O�x�H�_�EQ����Z�NVl�����]���u}C6��hQ�aD�tC�
ACk(KSk�-XN��P�X%8����ǖ��ƕ%D)d��ʶ
|�2�痒"�),`��E>n���&M6��y�!wWm����=T٨߽����(ё}�C��z����^��5��w,����F��^�
��s����j.
�J��D�٥�f�=&���!{���h�4�`��^���#V��.\��H�h��dB 2�V�'l)�i='���sm�� �5HK�4�@.oe`���m�o肧9��r�R��3�qK6�mŖL�;�����I�r�<˶Q�t���F�����*79HyUU���嘝��F�A�'��Wԥ��i�`9}kK�_E���$D3K��|gbb��$�;H�⑈"66��_�پ���"6ddd�}���� :7�)�	�diPto�+����<��2��;�J�
�Z�!����zC;5$/������~4�}��?�/KCK/��;_�u𔑬0��U����5���(�����{F@$u'5������#��86�sGl>��7����qz.X�W5�B�vxH�tA��à�Ya&i_���t�7���5�l6�yÓ�<�v�z�0ӆ���:���ۻ@��P/! @��8L./f�u;��ʂ��Φ)4���������mRfd���:p߭�^;<|�V�b������\��O���������� upʌuf�yVC��[�5
�#J��(ɍW>o���~!�<<�) Y�<���S{ֈ�����W'�2�P�K�w@ɺ������Gk��2..�YJ���Dj(�>!aw3P�&��^�.#L_Зڜ	"�����GrS�O,�D���H�J���x��-7��#�;7==�S����P���uC:��=Bxt.�%qɽRD@�{VzG�3���n�U�����0���?;���ǘ��PĴ�;�k�{"��_�=�P�걨,��<e�B��H*p�#��0�&7ϧ''c|���k)����И�w�����閉��-��H(ѝ��j�*O�9�l���sC}��Y>ŝ��2�P� ��Eo�X��,�w�Ar\	Ǩ��n�P��n�����#�{'�q�i
x�"�kw���Po9Ц�;w�p�C�h3�(��}����ZL۽="p��>�u��ֹt�Q���o�[X���=6�]���X�[vYC�usL��L#Ξ���<I�;A<�<�Ȋ��A.-�K�C���L��Ծ/r�1���lz_�����ϟ���>T��K�7z��qH|����"ןZ��JJ��U ��JHg��}V6�����֩{�S@m����{[�l�!�lP��PQ1sV�ꈀg�z��gB��Tb�a݈�n�����Qc��S(f��8���RH� ��%��G�zL4� ��篁� �J�<�;���좦�ݷ���]�Aev)�CC����</�����W���'''9(V����O,U�ʝ�"�W�ܖ((�Ѹ�:=gaa�?��:6��sZ�zX1ݝ�{��o����Q�YQ� ����Y�4�B-@�.���rP��OF��L�E{2��+�	B:�. ����2��6f��L��z=�>I��,I�~��=8a #�ũ,�}fu��Qir񰶾��ݻ����+.w�?��o���:��G��Ȉo'�.�a�d�%�T� ��T�`kKg\�+^����)E���ghXL�g"mȐhHw��7o����w��[��LMɖ�>${'���U"*�x�����K��9<:��)���m;+���(��)i��p�����(��M�f�>ًv�xs���H�!��`f�`F�E��\U��>�--v4obz,���w�I�����Ñc������p���{�(J�c��G���-}C�[\m�Z��f��H-�[I�"�gf�il�>V��uϰ�Bs�33X�RsS�!Ob����gi�N\\��c��b8:���ݔ=����͹5�6O-�8$���/�cьw/������<�KNa{X�-��8�s%h �Z���E*b�>�b-h�R�W�*�fd+�g�H���n���G���H��������|t��!��5L4�B���dRVT�W�KZ<��a1�4� Ղ��<��@R-��b��(�g�|��</�fo_̯������o�wx���7���Ŝ��}� {���K�ȧP�a�H���A������]02�
��˶�R� ~Ä���9.���F�d<�q�) ~�;�DJ>"t��lc�G�Y�o������1�@�
������?I�T		������{����mݷZi������f���	��p��
!!!�z(Ԇ�~~��o��G8J��4����q���D�%<����L*f�r�8������&�����v�5��iL�y��W�)�F^b@|����z�7HMҩ��W�Z;<�j�`�%~s]��{���Jc������.��c4BG�ȿE�k_*Xw�J2.6Is|�k�؋<�3-��̎.�]ў��v�����.>����ohBh�k�[Y�<%FtE��3��{�CJg��Ԃ���o��ǫ�+�؟�y�AtW �F����M|^ޙ��SS7��#��Ǿ��� v#3����Kߖ#���2��^&�%����^�2k�>!��`r�Y2����i�������[U$92X%�\�j
ME@���80�kWHX��W&��kݽ�¼��_ī�d��Ū��B"Y$Ϊ���d8��AE?�'�X��"�,�~��goo�4�#��),	�����M��}��<o��Ѕ�/i_��YL�����.3iQ��z6xǨ���?��-5ukx�d�XNN��'Hp>=l�ސvp �,xm���>(��e��f��d8�PYu���c�6�x�:R��y7}��±E ���������נ�5k�ڋ�ZE�p�=���Q�,��8���p���1U�YJ͌�L����w3�PbW�����k��«ޕ�\�h&����O�&�K����0b/t��o�QeiCYƮr��j��;��d���}�&��u��7�^�iq�o���,�)���_N������g�E_��W�b�$�I��ژ��m���&S��|I�uX��l���� \YˬB���]r�!7<�D��ǊL��(T�~��[��Ɛ�ɵ��(�&���S�J�nn����o��>�{�:-���U~{�ny�^������m�XTT���/��Sy4:���Ξi*�=,�^<�:/���'�H�������6��ϮAv;��?�0ߨ�.go�yV4V�|%��x����}q1��-A��@����bח��ß��,h�J����뇷���kƏ�a8@��2H~�(U蓪[�-0�=�H��!�������Œj�-52��Q�`��[��Xpz��F��v�6Y�
�6�ф��,[O�g���i��B%^����-�N��wBd����X��y�<�wW�� {V��nDV麘m�q�5nM�Ϧ-Z�$����s�<⑨V�6O�%9jr&P�&ED�7.�VWq�"��G�gml�@m���ojo����b�:�FB����ԁ>{��'����o�*�(m�K4!�q���d�+ό��>�7�~��9f�^Y�P�?g1`�Xg�% ���߲5TL�-s�9�E*��rx�Z�LTJ��7���%:ߙ��%J�}y�`q��u�kSS2&�|?�l������
J�ͽӥ��5�z
`���`�:6>5, Zξ<���PN"��(�g��Y╹6ä�C����&P�\�&�,�'&&-��#3;�
�G�rF8^_�O�V����^��=�X֥k�dC5|@5��g�EPU`�~�p����6�~���D��m-����F����j	/�DK�Y�kd�l��QV�gy��T�*w����Y�~-g��Li'(�E��U�Ը6<�ss���������U�w�
/dM٫�5�M+�/�?z�.�t������3j �]E����^�N[���d���!��\�.������&�+22��a�V��"־o��'>�a��D�<`M���cA�&?�I�-���jH�Iy��A1��0��,)��mSH��J�/���<b��Ukb�(<���~��̷�w�xw���`9:l���1hWFmʡs:05���׵e6tlll�&R�D ��[�H�Dr���V���F�����ӄ�.���Mhg��PR��?L�e#���Pj����{�j�e-�b��V�������3��1��'�
9���=���\����A��[PDw�4�$���ݼu~��i��my>��͙1�~),/SoH�.h���tf��� S�
��s���b�(יl4��$%T�Ы9�Ǹ�@���G�x`fַ�C:��Wmk�½4����S��|�K��/g������!�X6s����L�
C���Iy��naӢu�	���p����ŰB�~n��PH��dU�g�5&[����?�2jy����6V� �_S�9�&��&Jt�v��Hb���C�f����V�C�>j����p��"��/҅sD�޻kY'�19LH)_�}������bJ;\�]"g���-��j�]���!KYYni���]d*n���c�(�w�����-˿}���nm��K��E ���Rq�y���}j*=��{}P��] ����Ĳ��û�s<6Nf����[��E��-Ȟ�e����R&�H�%�}���>̀ ���c�N�޻���[Yy�ߦF"�@$���1^Q���wf{l��zy�Z�	�N��2cj�~�%�r��Llu..~Cذa��=@�:CE�M���ٸuJ���[y�!�`��+�|^NN����aY��Þ�cçD-�V��w�� �}(렙@Y����Z�ų����u�v"��u��->�gu���
dj?�ɉ����r��9ƞ���~���[T$���zà�(��S_��tsy�n�7D��q����o9�����T�>����Pr@���X1ȆN�E��0���M�PyJ���_��p������/�ܭ�P����IrR/c;��09$c*�&��w���)�Ԗ�('%>ж������{�������\��:F��[�r7�$�P��o�/���O��9 W\̝2�y�U�Q;�x�j�nP:J�IH,�`��/T=^�wp��uμJt�D��
�������{<R-$j��*�*����,�*b��N�B�������HYh3z ֐��)�ƵϤ h5�����A��Ik�Q����e0�3���(�""8$�I���1�����I���O&������s��힟/="
���}�����d��'��&��2�3G�f�0����s;�ԉ�"
2�4�ƀ���Tt�K0����1S�1qҍ�=��r�Łv)���O>����&��66V���C�e�nP7gޕb^�	�'���J���IDF�fs83ֿ�x�&�7d�W���~3Y᧞�=��n�('}S�f�h�	7<�Ƭۈ��H�P�gx�c�Y}_�j֜]�(����cA2"pp}%��͔12����
ä���d{q����HT"]*���[N���w@r����1st���[���NJ��㶵���w�(�O�A�:?��U6N� ��|Tc�S zǈ�|�J�!Y�zidA�[9����.�:��i����C���!a� ��b���^���=k�nQ{������J�s
Yḵ����8Vm93�P��{���"�s�wN]���)I����������6I�x������*�r)���&���ܜQ�����ty�j�`m�#����9��/}��NO�+�]��/q��7,/��v!�v?��Ս�%���vpP�����\@�x/
�Q쳖�z��*�Ez�* ��YX�F�d�ۀg�E#-,0<,�030w����a�,!�}\I�4ᵶz�Ū�`�Vʉ������bh$�О�
�_Y�42������+�q&�i(����_Mv�9(�F����mU��}Ͱ���ۃ�G���V(m�ti��� P��!h\�:IojlD:]0~!E���:n�N�a�����I������8�z�A���>��#�������c�%ķ�����_�m]�}����p�;!�f�#S�u`:f	�����$�Ps'������د��F~b�a|�-��Qm5[j)/�p㖿�Hc4`Y3�1���F�iio6d�~����M!��l�-��s�}9���c3́%Aei�Q������5Z�a�ݯ�㥩*���S��SSߪB���24�G�r_�[jk���I�dƠ��"2��1���{���n�'��|�Y�MSG��jo==6@J���Sc�M��7f:���MG)�B�v��a�Z�K���׺�z�q)X�`�`�1�-[6��o���=�Z�+ s3Z\�rKOO�_2eF_Ǿ�;��G���O�.�"��Ǌ�a�,�s���*[ ;��j���|��4uv���D���4�q01$�O��xđ0+oi�r�%�|vky�b�����sZ�:����}����KY^lH|�6��&&��`�FCTl,��g�����YC���zC]�$�y�Q���l�����-��H�u���`U�����+�����o�4"��6@�������k@��$M�}.�����]=�z���𜵵G�=�R��2��Q��B��[ e_XJ�bAcctoo5`qqE璌�"�����G�u�<O����HP��d�.���g�mlp�rßqS.�_qy��p��l��ݻw��-
u�k蘍��oP����۰�����L���I���F��� ��1������CX9�~�xP6�B9tSJ��i��rI&�l�6Ǣ��>�4>��O@MQ�AsRs�u���8�8�s3O�
�{�=������Z����w�� [�ҴGɮb���t8��_�<���C�����~�nm�e���z���Xq��@[�A�'50@4`ř��ϳ}���%���C����v�]�2,H�mo;y5r�남��9�ԝ��sQ��iV��'#�R�"�*����.��X��i-�AFjI?�z�o�ߙ����
l�J
w���5c�e��>�7��n B�Ʋ*Ԑ��U�{�J��/��{����BB��Ռl�%i�*�)zn���}�
�~]���ORj��(՜.Ob�L��}�^�]JpggHRJ�.��5�B;*���6"��p���9������U^���S�r��(��	4�"I��k�q�!q����bs~Y����)�B�6�xꀥ��C�u}`Q�'�m�0;�-� 8��]&�[�S��P�x�nR�{��:�� d�Ø���)n�ܸrK�0�o���ss�6s����;�s����C��h�W��0Y�QbvvQ��ႉ��k)iiHd���=�&}_?AB,;�"��8|�l�[ظ|��J D���|������-���9#uG��ffO^h5�;(
5��^�W�����Ĥ�P�N�k۳j5Rp���z?����;�� �6P.�s���5�-��8e�}����xJ?�ǁB��#�6�g\�q�!"b?+ ������S��x@����%/}n�M}a�9<��9���`�6���~X"3�iJ<�|D���������I��	K���읚𑍎���j�sߵ8�]]�Rɭ���X�]\\|���a ���$�넪��S��z��/(�jY��|��C�`s�����&؛E�����=A�D�*��}�"���ރf�v��%�:|����Q��QQ>��0 %��t��Hw�,��! )Hwww����,�%%�������+ҝ>s��s~���⸰3s�ꚙ���*��8�&�y��{�y��s\\O�6�������1����j�����e����0�x}�����*I�۞uNd�ሇ�w��W]�[���E�|�+Ra��G�iL����-�.S�1���:��8��+��:��������K�3����"/���+��}���^qo�~|��X�}NsɝڵYՈMz�mN�K�m�����tW�B���@H�c%��"n߾psY�qޙ�$GF��C���`��]n�wv���7@��
��Z�7jǿ�Dx���ׯoQO�-��[��� �R
�����1�p'L����ZZX��O/��r��5= �J|!�7�팋��+��_�� >~=�K�K]O�ymȞ�Z=��E~I��e���Q�7��ygg�s�7�888�E�q��u��}9��_��dC@D��*-M�<��0� X&�zC��jO�e�80��i2�����H�߮�#Uw)2�{b91V�c	��^ ՟rQ��*������Η_HT�Z�6�;��ݝӼo�;�v����o^w����PQ9a����(
�}wP1�T&�
+*j9n:,2� �RsfR|�
�W�O~��3鼕<�`i���`���KY���Ip����c��������Ze�����I/�V�z��WdB<�,�6��(̛�b�w
�����cE�	��1AЇ����:le�p�����TRq����F��跉ec�;�F�1��������o�b���Љ��m�f�D���Y�����ֹA��(����yN�|�53q�e>�͈�s:��iЋ�x�'������	WW������A���G�D�L`#Ƹ�(t�@x��S"�uV�+�����1��H��j�&�@F)Ϟ]��*�B�I�%;O=�H� �c�H�Nc3�|?x#>�75����	+�
�d!|�ǂ�����?���;R��r�E����,��g9x�hV~��002����5R�lU���2�C������� �C�:��ŷ�[�t��I�С"�\n>�`d����@Nl\��~=0��������70z���	�ۓڕ�/���mm��{Pcٿ�����&��\Rbj������6��G�b�� X;����m^dވ�y�ų%Z��cu#�d��x��v�M��������^���m�s���d�kJH��3Ux&��,{�~�=�����rdك�痡�@[�T@ۛ�.;j��9������趋}@��q���WH���ncj���t���"��vh-+k���-e*#��а�����?�XY|
�h�t~�� 
�"�����l�b1��"Ɨ6���f��m��%�\�U�ŵ�4HY��������u�5�t6a+��o�j��b�;����ȝB�X����'< C^��N�§������p�^����w������W��7	
B�t�<��w�~��_G����̜ǭrh.d������$b�#(�:��ũ�3������!�����:T�(rپzl�����؈T�U�MF���`GEv�����冷iS�s>z<ݥ���v�×�6����=Iu��do��K����h��P��y���hu�`0o*�kn"Z��Ǚ/���	������'ѹ�|v�wT[,�*%���5�"� ry
��>�(3 '&2m]]��p�vMLp�D6n}�R��k+zя=��r��xe"?-5u7`�����mͣE4j-����6�ijn��E�^	�U(��96�NL.`.Ҹs*!�c>ξ_�@H�-ͿΥ�rs������%555�D���k�{���]w�=�i��B�0FX�>D���f��hb�ͅzyLR�l�=���Y��p�'ė���Η�|�Cߵ��>�����Ed�ںF���Y�{Δ�,3�)����#�wAM����Z�Р���^��ii�z��������mA�I�I?���}��n�~F;�8�ba!�/���{�ϯ��x��v_�+�nb9��GD/�w�,~i��X;8(�N�hTUW{�����&�x�����|YȽ�w~?AP�%r�rE����б%�"1�ھ|���] *�1kZgD���~,OE�0�}�l��C�g����~V���=���&��N��hK�LhK�5�<��.u:��KD�HS��)�"��oW]�����4;�dI�|�R7U���z�֔�:$��dm���ǏX+��f�<��~���ܒ�e@ 9y���
 C�X�������_����� 4�y��dNd���u����{�۔���s?�-�A�����Ò��yv���������v���cz��O��fr���f����^K��k���)��2������$���p�Õ��4�IW^���W�	&	��7��g6$��­���]'��m*3${���//C斗�Bca�����>����Eo�l�P�|q�ւ5���:J, D�R��w]�u����ggPg�чJm��������8���)�ôFl$$��ղ�ˡ�Q"uMM�elXᅅ,�ĉ��}+}�C-�HA�qS��qHk���Ņev�� Y�3�bVNL��⼕Y�3+|�?��~52ӫȷ�{k�L��lJ���8Ą������_=I�x����0a[��.U�{3������\���-����PfH�H@SK���f|O�Fsy�h�FUMG��v�(������w2�|Y�!}�O<=�
�KQ����@꣓f�&"&~jn��Ǝ+MEU��w�d�$edꌴ��avT��@g��߀o(*%�|y 2F'FKCV������IDH�Ch�+�=����𹶨g�b���.Y��3��}��q�?M��|�u[�y>Ҋ����N��<�(���	����e�������,@4�
X��	
�:���ǣ"g�[������K�����XU�0Hs�'����x�,oim=�w۬s!�����'�/?� ���_��.��1��%�y�%)yiy_�e��aY5'������a+��:w�Wll,do�9Ҳbt�>�R� /���G�����/��L��$JJ˼���A�gV׮-�=��-��^�.����~�&�� k��K����7�r2q',���[F�'8&~�_V��[^�C�dk �|���e�Lg1���;�Gw)��v��"��9���==#��nWyHп�I��f?6����H*����)_&�������#��O��?AY�:���+~֘�vD�݊��O(�����)CCFĦ�'q�	�ܻ뉰\M�9o}����.�������)I��x\�n���];�(j#����U�R����Q,狭d���ֳ�������s�C���;��v˥F��8Cq���	:���DuWv��;ᨯM*0o/C⡧w��?��Ȅ�T]�U�	l�z��%��'���\\\���%UkDe�{��&�0ɩm @�#�ĩ�<JK>궎��i���S_��s���S�hδ��1�F��2+���dm��PVc�t�l^>���<	��C�È՛j����ن?*�����{p�-�9=�Gؚ�v��e��++lm��G"�YUĞ�Ƈ�6?�
u=:$a��
#�ĭV8�B�ry�C)$0�龮���`�����V;k}�o̪�����w9�R������lh�i 2i�ث{��*F�/.f��� S�P�
�w�y�V��b�[��������H4���.�y�H/$�3}+���k�30].����Ε�����נ]����{����z�8X����l`���tTҜ���3�b����%?���@��f)Xb����? �#���yh֪s����$��=э�[��~�`	dO����q���'�d1���Q"�=/�~����d�a���uT>�1��	 �9������:�Ur��;qp|l��	��--�^�f#�����[�hSp!˄�7�'�.|��hl:"X��fb��P���Z��&Gk����(�� Sf���
��-���g��d�!!1��1!~�����R��u�W��֞��1S�얠�t�M���d��M�Y�p$��Ry�#�"��j6�P;wF;"N�Q�&���`��.楫&�遊�m�#'#�9IB��fǖ��[��#�/!��QmR�=_�ɕ8<��R2��M%�Ð�lEmdf��n�9��#� �%L�/�!�ZŠ�7���e���$�Q��a��ddf�%  �������{����=_�I���I�x/�����8��3o�æL,6����+���
1YY��v��<y�����.��u�g�=v/���KXh('�ꪛ�fm������W{�#�mZ��阙'N ^�^0���o+�>A�p�q�/�62�Xh���WM��R;��:ڶ�Y�n����NM��@����Tѭג�,�~��Ti�}!z�`p}{-���9Osi��Xz�?Yii�{wщ��0S>�&5�D�ļ�"��?P�W�8ݥV�r�g=?<<4>��ZBp"�G�B(`d� $q�_9�@|z�I�v]�E�ynz�I����؜���ٜ�+��k�}
�!���Ǚ�0/0����m��6����`%���qP� #�B���4��� �0�<�	Bb�=�©��o���Q�0-�4�����>��7��M�ŉ/;����1���mϬ ��WI���o2>�q�K��ɪD[�o��������d}����݌�JLL,i�@���'޵}�#�Y�������������zK|覫�����Eж��d'|%���)&\���dA�U�'�83a	;r5��Iʇ��Ȑ��1���lП*��rH�橵+�xP�bc���-��ٯ_�y����wŷ���>7�61<���h=�J�������� �dȨ�ػ�3���?� �>��Y�~�CL/�a�$N�|�i7V���GE��SS�����#�ohj�C��Q2cA��J\�Ѯ��']Y���w"��L��eX��=*E����/��*%��͝�����˗���|����-,��#����^1�mE�>�"��@|Q{h���#@�>h���.)-+�7��|����0o4bO�y__��49S�t�&(����
2'������QT}�� G�_���eI�������J��o��۫���.1>\nmͰ��mE;���;=]���!}�)�1{vХ2�k��~���pC�����O�:�}_On��V�'H@Q�jAs��9t��B��Ԉ�O���_���������"��>^��a��_����e��z�
oi�v�R�rM�VM0��*�kYOwoo��svZ��:����9A����#g��r�VV�,�?�Rc�Gs&(��`T��?��J�Лiq��tO��}�����Vi�y͆m��-t��Z��PR2v�z^��k?{F|��DDB� N���+�� =}���7�,����o�Y��Mo�R�~_��_׻�~��8�`�!/�z����OS���2��<5�3��8��z�$�ܰR��9{i��Ü�2�a�gK����d�6��Z�Q�Q�UGp+�#$Kޞ�.�e�Ff!Q�zr�A�����j����1/��S��ՕQ+_&fv��NXNe�8��$u����#�Y�P5���^����>�<Ɂ.n4sQ�,1�rRXC��:�cbrA���^�Cvp`��;9_&��9P�}��;y�Ԅ/���,�#5�w?8<���p����%���~]ږ�_?�h�IB�`b��e��i5=�'�
O��k6rݫ��翺��5ƌ�49?�｜<��^$"���$�Ǐ_]�Al~w��Z��-B�1|� G>��>�&\����^�'�6h������Z_�*o�/#�7�����0VU�D ��O���,��S|d�ӗ�-��w�EA �PRQy���l���+���Z�ww=�[%2�G`��@���$�#�͆��{�1f�jv����σ� f���l��	��8h~�������W���5`他B��I��O��i�����!����=��L���(��v�Ŕ�/ŃMe�_�.	�JW_����:.ٔ�
�wk���׊�S�JEEȇ���u�u?��ؑ��.�{�K�/��"�&!'�;z�X:e9�j�����
��+<�IAaa�*������i11�*I�a/��-�ϭ��;��t�ﭜ���t��j�s*WCg��*C��x��X���Fv�����XV�16��[o�_]�4��Q���Ȓ:����_o�q���-�utxx�EL�y��[ޡ��۶���ᘥ�/ֽnv���P�w����5������^��2w:��H�4����(zt��A*#����iq�>yW��n���%���/!�����P��v��3_���jW�S�|k{RGmʷ���OA�tR���d�UU�� O�Y��_�nRi�?$b��ikߌ'��g�V��辽L��MD�O��N��qS9����U�[���k�f�پi.��y��<3�Wq&O��\ڷBo�UL���[<8B'��s��-Б#o��X<̶n�t;˻����FG
0z*��k���X8ן�����0a���Ne�iAp���i�g�k�uz?�\�D����z���Ȓ;s�X~������h)������[N7�	!�2�3��ٔG��u�K��+5��۴_"�����|q��'Yn#cq��h���9�&�<��۶,�r�_��`Z�c��e}��~oo{�o]c�g��Ǥ�'�09�-��_�XA����;��q�����C�����.C������#�i�_�n$§h	q�x��N�Y�C��ε�U
�5�-&�C��o%fd��+���95t�,���C��NEm/�>���}��ݺӆㇶ	�`Fj�ɺ��8�Z;Z:|캖�,��܁U���T�Z:�K�1tOmO�GJ�^ּ�v�6ō,��5:\�g7�;�T�/�e�++��]`t)*SssV�k��X�}���Ԅ;��	�4�T^^^Ō���II^�*��-c��"@��ו�M��,0d�3���42d)T��vy��F��)?��S.8���8�v�iX
�|u�m�ǚ�ƭ��C�*�-πmQ���p=�u���}��N�}���l�X�߿��<��yI���Q`������pcjB\�㭠�B�I�+�Ծ(���ۆ�&����ɐ�}�'㵡Q�����SW�%/��;����umE��m��^8�8Lͅ��(q�mk����N�.��4���ɉ���Ӗ��[�LII�۷�i
�x�^�gO�L�M�;���7]$�w{%�GPay�v�S���F���I02��@O�.�X�Q�#E�[m���r��\OuUA�����Ɗ��������4ˁ�U*/���bk=�]�sPz6��io/Q�:���R����8;�#"Y�_�6T'W�E�?$Ŷzpr4��p��ZTzv����un��G�v�򜁞!$�$�"st����3�4)b�#��XI>��&�����=�dqi���������P�{(Ԉ���Ü�5%fR��~��$Ԧڋ���{,$9�s⯢'7V��aK�_ZKfƟ�9ã,LpP�Z��\��Ɯ����&/ػ����B��OW��n�UVpwK�&�a�ݽ{7�R��%Tij�ǃL��1�Lx��+MIONL�&��|I�-�v^n۾�:��Q,'z:ha��2K�S_(�sm�%]4b��Ҵ�����\�@�s!us3�������J�&� ��ޖBG{K9k}��VAߊ��x2�8���>�S��!1��XS>'�}+W���\;�
ޏm5d�{���(z�1�9� 
���@�<gG��e�9��L�8�%��$��#�k5ߓ+6�aJ�[:<���		z�& +Re�� {�W虘4H�X:9��L�{��RUe�y��-�Ք�����\��d�,��l6wv�����H8f'���wp꒻@��Pe��@YdH��)M����|�(��J<
���(�0�ş���*LJV��jr�uVzw L[��o���
(�Qm�m⢃���l�]�e�ӝ(��n>p<4�ʻ���N��C8r}j�>�Aqn���a��g�՛�@�� ���%w���pVn����1������n利�?M���+�sU�PF�9�df�M)4��S�J���ȽŴ%6d� >�y���y�V#C8�.�%`�ݥ�&vf��ꠧ�LFkA;q��������MϠ1�n����3l+�\��-!yj�cx`�ɒt$�����DCs�� ������
ۼ�VRߊ`�Vn~�J)�=��z �''|��P��'�zm.���އ�'r	�$�k��/Eғ�i��|��Ԛ5@M�s��Y�i��=[lZ����(�_���㝜�N���i�Q��^c9�8�>X�9Ig�j�uQ4yP�$
j�ZX������z�$�yz��p<�o7�X�����+��kE����Bs��S����\+o��#�Ѕ������gdİ������軷� G$��Vu��x���d3���4�6%&����B��oL��$B��!��R�:az� L`�l�q�L�8��gr|�a"����B�	}����or���Ń�^��E%Q>UJ�2gء�]+9�C�����!���OdI��^��������B�q�x~�S�����]g���9W��W�Č3 vAdr�9�~�(CX2 ��[�x��9��0_`�:�J(mT�Alָ���xr?�gkce�)W���Q���n��Ut��ɟ-���$���p�Z�_C�w ~-8{���ϥ8W��7�(�Zh]�5h��s��u�6L�����ʍo�6���^QR�ԭ�����W�r��L���$ʏ)*")�|���911T:�v��n>mǈ!AO�1`��oN������H$^ٯ�DLJJʝ��L����X9�`*���-.�[�q���a��`�m��i�
�c�?�*����/��D����6�ʰ���qF]]��#�W�|t$�oФؘw�Vr�HijI���v�{K��O9h�����6�&K�k��o_�npa�d�I4��j.���y�)�AoR]�Ph�݃^BيY�g�������=�S^.���&.���(S��{�u�l�w޵�E}z�F��ٲ�k�N텳�����Z�w7��,�7��$Y\$nT%�3�����	rG��wg:ն�����ǹ���5^R�2`T���ٿ˹�Gq�.\d�W/������,��Y'	����(�����|��f#���($�+z��I'���=c��|����s0��	nE����1�C� t��ȓ����r%�@���E��qKܜLK\���C�y**a�����U��/nmz�>,�Cz���k���Y[_�w�x� ����15qJ���5 ]7���O��.�껺bT)B��Nl.Ϻ�E�HYY�t(���;/Vk�c]�K�3�.��:��M�[,(�?��p���[h�9�HT)22���e``�r݆��?��+>wp� z}X����iq�^}ش��h^� �×� )�j��s���X�X���"�]74r����m�T�=X"���ź�O�����m�g�������C,x�k�\��$����Ms�h�ۂ���t��ܰ�[c�PL9<�65?ˌpL��b��o�	#╿�ʹ�a��E?;��)�,;Ҟ����2 `���#t	6�XUB�r�|���e�v�h���JQ���Z/��+��
A2J�����,�{� A�!_k�աuw����T�C�_b**�^I�$�����m��a��E}�D��ׇ�R��8P��pvu���C�5`�4P"y�'�+��A2�?<%�iI����Y��Q'h^�7�<��gfEX����C8׽�2}>ޡ��ʑj�Z'�ӑ�]��v!
m��f��^V9�����F��M_��{/���� R�lRbE0�\���R��^$ҵy��N��67���罽��L
��ϻ������뻏�b��W��B��N�sv>�z��-�5��vQ��ܹz�C�׮��"黦&�)wz��%��Y�@�)렐��8�
�>A�LgX�$~���~�s�}ޤ�ö�~���/o��U�s�r����T�#֒�l�JTc�	�����'�*��k�J|.����G����Ax~I�n�m�׽��u���OU��@���3���t��u]�G�<ԝu�Ŗ�{�;b�p)ǭ���ۢ�Ti:3���� �����]r��+���xxT�C�s4�Ss$�K(�8A�ڳgĜ3{0T��S�v���))�KF����N;<In/� �9h�(~��ߠ%FdA�\'GM(g��|/0��	�Y�5�7�f����n�����Y�)eQ�.����+ƪ7\�ZZpl��We�a�)���� ri��|!���h���/�����T&y�v�z!�O���&ݟ`������32�U_�Sg�;�cc�X�I��x���P��E�����mY��$������3*�5���`��J<��T�W�� G�Ǳ�h�_�n;!ȌYҍ���tTJ���D׎t�UNn4��ކ߭��
���ӹ�y��;������o�h����ᑥ����P�B*;�(�����n\o%֡ #|V`��t�=rӗw�9�i�V$8�yT'�YJ>�יN3
��&���\z���؍���\�5��X�Y���V��(�܈���̥%�q�">6iO�EjkZxE�}�q�L��P�ߢC�5M ��L���-s�	��<M��4cJ���˧�T�=?=�ssݵW�n�ߜ���E��n�<���[�k0��a���^�4+P\��jhz�Ʊ)��R5vG��PϽ�s|T��[�����vy�Q�Y����;�+~�)Cs&��7�g?/q���N�O6l�<�̚�3hmmc�s`�Ά���X� �L�S�G&œ��o�ί}Y��I.������\p��"����ܦ�
.�vh2��`��=�$�D��}͠rV��B���� G�HD�ƞl^�7��
Z���������@�v��'u_6~If���u�M���Ǔ0�=�dk�?AFGd��qm��������"�ڥ�5r ��ÛLهa�**$d�C��V4,_>�]��p�=��-��lNY(+�-	�֝���6f|6e�����;G�|�{��٧���?�~�ntӷH���ō�l��O�,���)u���M&�%ni��$#$ͳ�b*O�[9^����v3!�B�:~�g^d0B�~���ntX'p%�MJֹ��W$z�$�w.��l���$��� ��@��I�Xr��u�L����i�����X櫻D��.�\�Y<`�Bt������.v/����Y
w+�J�}��jK��X��������hv��E}%��2�|*l���Y�1��ϯ]nj���b�u!�ܑ�ud����:1L�����.w[@ظQ��&��#E6���������3z���=� %�i3C�%f�x\n���b n?�/s0�����~��#k�C�+͋Py ��M�X5ĳt)�/����.��g,y�h�5�/�TV����9J�~-���J%
o`�ja�H��J��2��%߷�ɒ���>��o�����*ྥ�s7���)���c?��h)�,ʺ),1�f�3i@NS���o��-�/n��*���}dJ�F&ff�P�&���F��4���z]�Xk������g����v�q�l��߿k��;�%�^�q��CvlR���B��O��*&���UZ+����ţ��Q�j�2��2�u���@�3����Vp��Yy�"�`��}�]���)V7�ѻx��\�]����7�Z��*�P�X{x�0��]�I�W�B��W��-��CMY
(�_��茸W�a��� �0��ܵqȒ���m(�v���F���d��<^9	��9��Q�8�v���RҤ�wM����b�����㋶�Q���;�7�}
���=Ʋ��y�j��������4�A���{` ��\�����x4p���hϖ�'u�V�0--�,��»öךLƹ`�"�����y�:]QP~�V�P����p�l�X��l�a�=�*y�C��>um��Ζ�C7.��m)��7
T�N8�cI�9�n�_i@�!s����\�k��m.
��Xx2�@�k�I��U�O+�ٽ��X�cmӕ��5��o}s�og��Fw����R�C��#u��*�[�������C�]���B�#��֓�%��RN�^Z��я���Ε��x��qNw����>��UW�|0�=)�/xc�ơZ���ܵ�b6��\'h3��I�k�!$�����V^��~��
c�������j��Q>��M�И����cn"���a�Rd��✌B��
��Up�jR}��E%��Q%��ݠY���h򾿌霬R��p��}
e�0
����Q�L���%(���^{�_(�$ƈO���r���7 �g��`g� ���;��l��	�z���><�߂-Mm�D�և�NIyyħOr�s_)<��qQ>~��C��s��K��Ӌ���˼���au\w�$��� D�vs���8g����b{�D�!x߁�z��q�u���sr|>c�|���0�2 ��ԕ3V��:�ȿ������D�,�I+�n��Y��q�bہ�9>�;w�|_�7}��J�4����Uw	���(������R)JQ&_ �K�D�&ZN������2��h�P|\���	����g�2�� �����|
��_a1�͋�9�cu~���Ô���tR�=� �ߺ#�2��;҂2R���ߧ�V���f<�r>q� ���"� O��ռ=���lg	c�u^e���x��q����K�(E��XAPh�mw��o^G���.��\ܫw�fܳ�1x��G���������lpmN�"ҡ��U{af�������/��4�*^��q��K� _����5/�w@� ���`E` ���f���z �/3 -��4RB�����'論��7����v�Ɗi0f�uD|�{#����L�R��S����~on��x����2''����3�X�"'�dnb�=Z�u���\Hjh���ၗP!%%%�u�8���<����rU�4Zn�y�2WT�������P�����1'�Bnw��U�/�P��]���wA��|����:K�w��YYo ��6��/��mKY3.x

�\F�w���>��K����v�s+$m6�WR�l�A����ÈF����EP�(g�ZSdʷ��,~��3Ǧ'��F\����B@�?��<� HJ��F�돕]R8����&RL��Ǐ��4���USP�M���� �
=���F(&%����Ħo]þ�g�==��T�%��G{J�O͇>5�/ېZy:�0��[�n�ZZE���6qxH���r>�����"�g�6$��ʒ#+.�Ύ.p�>"��
Q���N��xk�}�f|;��(�d�����f|m�[`�3�?��%�GքMu~{�  
P�'��Ts�7.Ed���{�#�hZ��L�X�Dd>P)�E(`��#�H�gc��|���)��3�_��	��Wt�Zt�q\�I�bt�m����W�57���)l�U*�ck���d�!�zR["(�?���t��Y���7"9���~10��A���6�ε�ol���u��.Ri��+��_ �r����E�6�K⦣��ra�z����:*�wӍ�	Pŏ����:��;g�{����qH�t��\k,�_��q��a����'C�I�ꔷ�����ɖ�����#���s59I�x�r���c&��c�ǒa�'����L��	�vG�5w	f���[�X��?���@��X	�c�'�N���5�c_һ�̿]P�:��Ԅ�(�`o�u���1���A�M���d�˰ 
C�6egu�1		Hbے�vd®��� m�mw�y��1��JA��ً|��U��;���g��je+7���Fʙ�)�9>���(�u
egWW������?<�o4��t`�3Ԫ
Ş	�m�G>������z����B���ҭ<�a:��c�{0l���'V,rG>�黑w��0Nɿ�V����sJ[�Pr˻�6ƌt+�R�Ԅ����Bw7}o�e�z��[`R �m���M��e{�0	#x.r�^���*�O�O�d60���XPrz�"��J��X?��j���¨�������܂��0��@�֯.�`�P��ɚ�Yɖ˺���� z�,���#̑��Y�4��թQ��T�E��Ǐ?|ot�\�^Y)���U�շ~��8v�/��*�?��*EH��_�SJ����p.\�� W����z�5�N���fM�B��TOȅy�����*^{X�0�*>�+\!w4 )u�.���2d�J��IkY��8]��[��a����9������:_"+V�Z��/��O^/~���F&&�?���S�rk�*��L���VMa2 ���l���W���{�Ϻ|:B�c� ��F��EG��܈ݭ��?Fڋ�RC\l������3[2�OL|4u`1<�uj�e�/N��w(�E��Ӧ<�q��`Gw����͔�3�]r�I-���F���-�j�E:�IH��7.�82E]��_��V�"��*��]�9��qǞ�C�}@�tTY��Wj��qQ��U8�7�j	�a*!OW cj��<����|�aƗyi5�B���SU*/vBԏca������� 2lԄs��P������\��"}��H�--�m��J�;g%�d&��z���RV<[8NB�4f�q3VE���fd>"�X�YoLL���]��,���g��ơ��y?O��<�v�8���⨾��=����BO{�z����b9+V�fi�>7���cô6�-�H9)��(��ˮu��	6BOO,������7��`f�?ִ2�\�R8�`�a%�S����z��A��>'�M��.�G@?\F�d����)=�r�Ț�GJZ���M�|��cJ�}����ɐ#ױ��w�\�7���Y�sؤ(A p�ж�x�ח������S�eu�+}��p��LǊ�u�=�%�J\1�"���e�"wp����@<���נMbݳ���+�Ş$"��u����59U��"K�hm.�u|���?�yp����Oѿ�ĝs�#�M��䶅"��5kkS>q>�A��z�=v�Q7TǦэC�!��PC������i����:�60S��Hg���&7
QVd��u�M?����\#*]�������e��G�ܨ�y�qF�V8�W"�J2�����m<ϙ�A������P�xlL���nN��ߝ���KYQB��`0�ϕ�j�Rh�3̝Dh��O�GSc�T�im?�8p������S>���"qu�W��KAW������4X����611Ah]?}C������#���q:�$��>H�'�)�l���'�q��o�]b�n��W)V�S�9� ��-�CFo�z<�׿&X�����ǔNb9FFF��v����`Ry��C++YhS�4�xpejSP��P���C�g�����PgD1��i�_�P6��e���8n'��9����A�8���Pצ/�{k�y�^���o_<�]�.�0Ƹ9�����
�S��cɺ<W��C/}��s�ڤ/�`i���hjiM/^b���~������%�.Q6&� $�XrO�/Kz��Ǚ�ȧ�S�pf�{�-q�P!��j���Ȳ"�Z��u�j9�2�q��Gtx��F��ň�Y��k^Vx0���n$Ϲ���0ie��J�����o����7�Dn��r�D~� ��Z�~�!E�"u3j�P؂�$���,��}rl�ϝ���sQRW��I� 3�x��lh
	qwCJp�V�#1@���a�@5���M6����kfƫ�֍��P�k�LQ( ᥽�!'�V2`�T#�Bp1�o�i̥����gBw6e���(=C�;��B{���Y��!!	�|
� M���M���Ǿ��,�8D0ӈ�&���52��(Ħ��O��]MM�V����A��V ��^svI��T>yv)��W�[�Ī��ƣ�9)����]ϔ���KƏ�� O)�>+{/f�mDh�$�YiSh{���>̹�̐$Tt�]mh�0��]��z�֯C�X%bYx?���o[��XRh'Ij�u+��x�aִhv���V���:P
BY��܂"��ɗָGOw��J��w^fx�G��Ϋ���g��vL���d��jYV�Rr����.p⸩逾��x]+���+N���l�s��r�pffF(o����Dي���X��;K��d� ``����K z�j6���U�F�(Hu=����<�"�����DZ�M�Y��<�ҵh���_)=1g���5Xq�L����b��0'�pF��������=h�u���%�ܤ !j��B�sleEJ�a}[���{�Ն7.CG"�; ���i�O�ho`���-�
E~"�	�[�����Z�|80%SSS�Dh����0�r�C{�H�����Z�x�_��'�Gސ����fU��ǀ}J��A��
.?�<b�1���ڇavӿq8��ЦXyZS�*���<oT]]��|2����/9�l���'?55Z��H�7������:f��F�����1�+1Lo��}92���������/�&n�IuF��p�o[���sb[��wޒ
no3qފ��K.�=�_��L��@ܥ�"����Rwr*� F�M���N���͕�C	Tht��9εtv��`ro=���ؘ��x����67g��3%¿{M�F����Ni���#6i��4��]~�˅ʀ��C�Μ� 5�D���Z����]������Y��u4ڎ�<@�ͤ��X��O��m��&& F�6T�̏�,�_���
'K���l FJ�J��m��[����!nD�������`��4(1h�	����S�pm���U�^�"& 1kkg1i�eKK���ץ���%����G�o�_��KDz�t+�T��*T%���Fd��3f$�N���=�G@@�n���=?���4 �&%9�\b��ƚג�����2õ����E�Z�0U�yV���#�
"N)7/��0i��2iiup����g�###�{�ȐǦC���bD@����(m`��bt��Ban�!
ms��bA_�豢(W�T���Utz�x���� ?W���x�~=�W��Y�F�����DT㼏�:��^��8>c<ܿ�a&L 귅r�LH�m(D9�n��F;6?V+�"J�,�ԏ�Ӹ
�fMS���hPRʧ��v"��Ԯ�5���X(��;
���\g/"���!@=l�Tm��,8@�4�~qd�����o�E �)�ou$�4��>-�{r��=���7���K�D$�5L`Rq a��Л��+�[��.X�5+''�kkv�6*�w�	� �x�_�<��}���gƒ ��c���'P�.���������}�ǉ�l'd�	yKƱ7���!;��{dfd��!;�^!N�N:���N�w��/}�����8�D�����㺯��19u����t�OO١���C_�,��ÿ��_�Q7������]�E�&m�F�[��Ũ r�/�ˋ�Z|,9�>gĿ�-�e�4�W�,x>ӟ7��lh|dV��A�m�la�d��7�'�D˃'�Z�dR���><�
$ �8jNDR���gk!�{ 
s��� ��
� �ݖ��6*�&?*��;3�n��.���"���V���B��7�t���T;ǡ�<ΠG���>��^�U��k-Df���w}/HD�'G��u�+���[_::.�t*��XYY�����[������G��,>#G��I|ެ�`vv�)Y�D����,jƴ� <���S���[�B��A*�Ss���;Q�{|q�%������G�\Q=������_�>�Hߩs���V�,��'x��f�3�u��Y��N-��،�y�VV�"�痟��Ӵy(;SUj&ydV��o�z���z��2&���2S� B�W+}��Sj�Nɫ����[}������i :��V�b�9#|�hK�ɢ8�ͭo�g�ҫ҂種�6�?�F�ڱ�]����"�W��l聙�L8�TU p��J])�64�����}5�>ԉR2�WK����߿/�8����L��yt��1�#(II��b97�\; �|���R��ɣ��{8�~�-��c��c	��3j��?�n���zn��4�'�=��<1���Jw:�>���~/��u���F:�%.p�M��X���6y�\7�Y�"��ņɨ�O����Uj���@�%i�]��Ij����LU��z�U������l��i�:�r��Kp�J�L�L���#e��/e������̥����E؏m) ���m2����'�8Z*u�Ļ���s��;i�P;�X���q��^_T��X��:L$iկ]Rvf���1$z�O�v��\~-�:9
���7��(ɱ��T0����w�8T�6��uͣ��˽Ġ&�ET9�����p��wehhg�u�[�wS��?�i�W��&�1�4K^��T��.s����HA�� ����v^:��u���v_Q#q^�`�R5���ܺeZg�]����A�NB��[���-��]��F�Q\�t�?-�lUW����M.��g2���_r�q�-e�ܭ`j/�k@�}�[EE��B?���N'~ GߺN����aݩ��]���ގ��n�rt]��SR�n���Y�?n���Ya�-a<pl�j�<���~� -�=�z�)p�,�<����ܹ�x/_�
�ͰT��~�2ުNZ9,��:]������M��;�t��A�\��Rǋc��3E��f�J)�P�A�?4��+�^j=�rA0k����"��Hw����r��
 �����סR�b��}�ʵ�U�Zet!��6D#b����4�XaY7�� h�[~R5 Ғ�+��gۤC;�_7J�����.�"��Fn��|�j�e��k\?�w� ���݊QW�|f ?[<�#�r��fQ���sM{i�$*К��+��q��)[A(�l�h�e�mp��Ղ�����
��_T	$�N��kԶצ������~�$����w�/����@�R�<�F���o$7ɡ^���#�ݹ��gN��g�+��x��]�h	H�Mh�޽�Bp�ɠm"Z�xԿ�BC ,���)�ٜ��a�*Nq��-��ޭ��>�>�@�D͢��$®���i�8� �2�klk�o���¤�+�.A��g�!��N�{�<M���(4Ӂ�?8Q����5�:0�*�S]�
�ϥۅ�vq{�����9�?-d��S}��r]8��I5 w6>�3q�k���sS��\��V��5�4utD���
9J�Z{x�-��n��k'"L��w�<�&\�U�bc R�M��;>��V�u޶O��t$���81�������*J4�4S��I���z���T��բc"��xi�k�W*���ꛘ�I�G�hX��'�2�=%����Q+uZEϭK�Y� �(~�jZv'����$�~�4Z	H"�jc�g��Tq/����1Q��O����Fv�P��o�X�x$7�,S2���Nς'g��w3�gO��?��wiR�����̧�m�=�e}���ݭ.>�K�}J]P�1e���j��n+R���f@}s�Ñ����b�h�������B^�d�<[鄋Y�x�=++%h���"z#�i����S�kO}�S�+��-2av��ٌ����U��LC���ƀ�|�_~��r#^ͮ~z�Ni/�0G!�>(J'���1��8W&
G5���)��ʱSCb��u��U^[K7�).�Jj��- _{��j���rpx!&e0��^��t�˝����C�����W���^ٖ�Y�2��C��YB�)H���h�n�i�8�����)��� ��{���:I�mq),Q.5X��ؘė893�,-wx�tB�� ��K��-e4dLu"?~XX��s��k~����trA#f��+���@�gty��}��F�ۻ)��Pé)���kJ�{5�zz�WV�	��ou���; ���H0����s��k2;�o�o\�9�QR�v�/1ʱ���d�U�	D	���<�ڵt����S:6
�R'���3���C8����[�uG� K���A,�60����(S+����,(��W�їՂ��N�7L��&�<@�5����g����ʃ�)�d��W���v������~��B~���jI���T@:m�G	<h���9*A�O?�oKY\�� ��b�Φ��� =������)�Ù6I�����wD�@���/H�J�^��as�Ȼ�au*A�6�Hŏ;r�w��e���-�+��:Fg������ϴ�����:�����n���Sf/pwK���du7��8�~E�,�%��Q�WW��Y�l���r�W��6ͽ�,�J%�DA�Q=�L�؉ّ�=�3�7Fr�'��a)�p�tZ�EQ$��굎 �����>햀�*��u���"0K�|05�<en�fG�*E�5q���D��^�;��/_��P�>+���m��u�aa���*`�}�ݿ��ktZ�Ŀ9��Gn�������<�7�(�>6��N�	����㱫o���î���^�*̍Ԁ'��9�窕��Kݜ!G��_�;�7��-"B����<:!+Z�F������z��s}��u�G�b��B���2Q	�h|��� ��.aP+�+�C>��V�k�+>_5�t��G!�f_������=$v��j_���-Kr,�R�XS��=,�jo�� �A��+Nt����m�%�K����Z���#�e�����W��}}��u�<{������"Ɩ�����v4� �9	�CCT���:!�߼����x��|6��"z��M����r����\���o;�`Z[���U���u-w�5u�СZ������Q�zu\L����ddG���u�@��|���R���
�j�D�5��g�91{k�/�al�b��U��=�\���[�ɿ`�=dV��cX�K:lO���Z�ë�\ę��yJF-F���c�J��KgQ�r�޽���|���"@���ڦ�U.��������>˗�|󩿜�\��Ȫ�$�(NN֔TK�I�������gF��94�S�,���*tp��aH� Óa��f%S����D���� � �z����T�>R�yc�H%P��2�x��ԥ<�GKKW�L�o΅UO����=|8zmٯ}���~���>����"5�>iT$?�=;�Ɨhk`�s3M#��荋�\_�߄g���w!���8�yQW�1@x
f�K%кs�H�M�,�L��0B�@���ƾz4���]V"[-������ZN��?��W��ϱ7��/v��Y�5]uB0�G�%uk��}����J#~�g�zb�P-�h�gVuf�Wu�˝����W��]-K�z���קD��Qi�U�*^��2MQwq�{�Y8��7	 Ua��)�Y���q�:ec��4y�xC����2�.�Wsg�o��p�w��<}ޢ����}_��~�]M/���ߗ�9 �;}����V���0B�Xڶ���Ȫ��%�Fuq�.#�ި:$�h�ͭ%��rm�v@���2h�BO.�Ǹ[cZ�J���c�+J��,���R4��z�x���Z�U���ܘ��Zgs�s��y���@,�����^�`�kT�7��*X#]�BK��5?��!��y�^�<��;��66�=�"9c����6�S�/�,xڣWˁ_Q@Y[XA��E�H�q�6��O�/�K���%&�k'
�� T�<}���}ꎺ��ܳԄ쩤�ī>��ծ���Sbb$/D�S\,W��s +-��C���tx�{q���0����B]]}Fp�ݥ�\�����A�����6%ԏ���5?�fs���ޣ��r��N�S�����slJN��+)+�c���S��7E�1ˡ�ë����pͳ�r糞�W����Z92{)��*��|�3k�4����NnI��*-Ӈ6A|�2�x���C�w�9t4 x��^�ZK�L�ۊ�n���BOu��x���cƝ>���K�j�&[$��9�g�$6@6r��_��R,R�/�)ȟu����I�-���r�!b�\����v9$4��u8��YK��x:�w����?�rc�������跡㝳r��=�d��LӞO.=�Tz������f�C�E7�����bDa�,��I2!E�yy�Zֳ�$���]����ZZ6�*D�Ti�)DpZn�M�Ն4���>[��g�35%%z�bE���_�D��X �/�.?����Oul�wG����V�b˴�Qg-^R2 a{���0�7x>����P�%8�]�.�}�TI�H�F��HFfze7H��JG����QL���7*��)x�6w���S)��h�Cn��4��u��/:w��ۖ~����,qz?|6�	"�/���:�?�"�9X�uָjo�j mjn����H=<T/�{�"89|��X���\�`N?&'�66o�^�����{rv���MC�etq�:4���8j*j������kJfU�t��d�+vv$����Q0�>7���)j�T���z��r8�'�=NX~@�ⳋ��C&�:ʥD�:՘Ca��e�ߞ����c
}33�@+{���S��찺��tߔ�u��O1]��I��0{/��Ƽ���ΰ���e�_c����'R�8�P��j���洬�&	�Q�`"H�ݯl`��~�A�t�����|,�N�9��r����
������_c.Rlu�/��JӪQQ�}K���{�'���$�����
_P�h��a�ro��}�>���N�CF|�B�� C��{���_�����{�DgM�J��jo�Y�i)|�R�������gi�"� �S�� ����~�פS.R.�8�nϗ�;}�pR�ډ]� �6��2��ӷ�}�"ovy[��e˃�lT0�I�UvAǎ6{3nx���meQ@���z|u�
$��C\���59#�\��V���v4��o���t~�XX*O�fu?x&֦�T �u����q��{U����5�	GZ1
v��Z������{?�[O�Z�O�Ԋ��WY�xO?�?K|��+�����쩼%��Ҥ:���L��Pvvvܛ�_�$����|�stp�����X;�4���&��SbB�bAsݕc�:H��%J��O�V /��S£�|Άhh��ܩ��Q�`��}A�&1�;�S�� ��n�{q�)֫����W���Gn��Ԯ�,�*
���<:!���&5���Ȣ"w�kL*�n?��l�'kN��b���	P+r��}���+G���T8iX|u���C����0^�W�mQ�ńK����Wj�K��_�S0(8{��;A������z�e?S�!���	�H�mmꗗH���xa��k�
$����a�O�S�n�G�ЖC�42�����
����vw;�Fo� SI{��Y*hȈ���4L$��s��6�����^?�ɯG�CC�nn�d���8F��� df�»��6��TӢ	h��3����WW|�V�M�2�h�
�0G�g�}v��7@�H�f8�ƒXu����5&�����~��0��pM������:�P�o8j�$_R�Z�ď�ٽ[߷C�>4����uCq�Ȣ�f��4?������P�ӷ&��4��� FKWs��~M� ��Q�$��ǔ�=�����w�3�Rq����(V}��������e�ݖ�DW7�����+���%��^�Q^p�u����� -b���`(҈�K0� S�q�b.��V<4^�m�5s����ݒ/B���R�܀7�}W|����f|��r'�8%��[�Q�xj��_���䚟����U7u+�����1V0���%zJ[z���Ŭ�������%���72V�R�1/�恊��h��*�X���{����7���ei-!�4x@`�0&��qSpg<�X�m���l_^^��:��)�m��Z�f�2� ��!�פJuA-��įr14���q� )A��'"�駏�X#j�f�[Yyx�\���������<�^{~�ͣ��^W�Y�Dy�O??;�6����H���WV���]��i.HO�������C�nğ�[ѿ��ܪn��#,ybb���x��� D��ښ�A�=]{F�D��A澎	��}2��~�S�4�d:<!��G߄×έwoO���QwZqTU)c?�L��J�kF�/����Vl���u��[�isb^�W[ٙ��tQ���xd����wԻ�c�~�-�SQ�W�4�^�yP�~|i�,�d����Ç��$�z�a��}?W�s��@�����������COKC�.8�(�����r;I2��G5����+i�_���СB��M�3��1�jC�-��T|�����<c��ub���hۆ��Yw���U8;\W���}BPv����>����O/cX�gi]�e%�r�
��TІ���_19��şs��EE����9:�����ܭӕ�Jc�0�ㄑsӐ�'Y����
"`^?���Z3�P��q�uڬ||���d���}�������B��~|�d�R�Y����K����)4ӹ0[�u��cʝ��rB�~�ܿM�&����ӈ>}{]��jGH�X��~<g���$N����p̱L�"^h\(r��.�>>�V��}����޿��i��  �Q"�������~!h'�E颔���? L'&|18�����K.ͽ*�H���m�3Ĕ��p+<?����Z|����͢J��8�4(^&��XI�'���n	�ɉ֫��e�v�HI��yJ]�j�9ƞ�^ljZLӀU��ivy�W��|���nbbr�5'��֯�L��a"��Vj����
|k �ۏaC�J�ll�����J��K��;�d*���Sr�
�|df]:�d:�t[Ƅ(^M��S�Q~Ƌ�%��x�3�K�_�d��Ƿ�?9eeK%���k�[ZOR$���ʮ`�z����ܣ�q�}��F mўA�*rZC��0$ �}S�t��=.��ĠN��5�O
X��W��ńI�=���7��i�ԃ���d<���3い ���w(ܸw�{�k������'Ζ��J%O�_?��e���P���N��'�Ǧ ���;���s��)�5Ga���*%��_��&�n�o]����@����Ss%~O�Þ`����0�5�`����}������*y�Z@Aǝ�z$\��h�hƞ�����H�\cˆ�ʵY�����=�f.�10�2==�h������h#�;������s�� W2ȉ ��gŌ�U��FʱӄP��3�����?N��{b8����h����"��:\���'���K���ޣ�ɡf� ��DS�
�T�L�8�˾������ʉ*��Z�ZUZzzay�8όh��aUX8{�C@h�\�/�KX��d�y��֡,�//��V
U`����k�ȽR�Oy,^W|\MD]gU4?Z ��ш���0?�B������!
�|�O�?�3����s����j[, ��,w�uTK��~T:�.,D:D��>��{3��x[WWW���]�Hp����+yw;M�MX���M�6�!v��������5�Gɴ�Z$0�Yv�j[��/V$2�G������ou+�Lk���
c:�`���wØŦ0���}�߹��R'�s9��y�dnJ,��a��fya�@����O�l`�H��w�:4���o���jL��d;�}tp�>�lf�L���MW;B�!&�=�٧��$&|�@�{�*ll<�Я�4���7Wwq��.p1u�����4vh�h��#x����R0�����?��i�:;_r�>���;>~atp��*Ū�B���/+�,����,��\�Ƅ>.�T�:7���y��E�g��J:������^*j�����V�d�ĳ"��8�4��ğb�w7�������1|�ňpwI*qx0��H4��mӅHfJݴ�h&�[�_��bۆR���7T:!ae�MM��GG��~���SY?��B"��]NE�	Q� kz�g{yn�x�)��uV�:�YYE
�����'_�$�'����o������J�0KQC��S��'�ŭ�'~WcS���K��q��r�Bu���x�:?02��7l[G��'P�`�=��&��ER`0�ջ�H#22���MS�;8;O��z6/�&cK�%r�˙׿����i���̅,���!R�4��� }K;���`�h����
�\� *mr�� �?�������J��!��r1 o�ӷܴ���_G�
8�o�u-|���KsB�D�	�ҹu��_��ς9Ec�d������b��jL�;O.��N?I���y����?=����n �]��r��$�g��g��z��Bv5jz�m��G�$��]�4��+�͋�z	�i�?r���7*������N/� ��T�ٹ��������z=����ٻW�|Y���#�	��O�5�x�c��3H�!�;B�v]�Qa����~�r�tx�K���}�:߸�E�np��3���iR�q�� J0Z�+o{�|.��35�O�SO�������22qn�Q-v@�:2I��i�����s��s����~�����Ch�=%�Wl��Ӿ������}���2=�?�u(�>1��k0�%L�O����;  ��z��F�P���j�����C�8�XHq{�>���3��qtU��Y8��+��+�A'��	��켼.m|WK�,yKJK��>Y�B�ዟ{�\� ��$�Ǎ-������7N	L��[�6K�`�;�Q��f2�6`	ع���v����A����t��a�/Hٱ��D=$ҧ�:�5���wP�8���̫�;�����|llF-Q���ǝ��C_��������6�.$OF����OQ,�u\����'�j�ܱKKW�mm�r��smv��2?H�w�t]�ʛ/�F�6�DC����?�z�iIu���"��Y(����/Q[��5��n���?ݔ/�H,qsbMg���u��Qৼ��-�(�ߥ���%7Imxq�{u]W��"T�������6�4uݧR!��Ζ�-saD:���/_��N����y�Ŀ��=4�S��|{��[X�Rb�/���C�����A�|'S��#���Pg�W�-mZ�U��AKO$�5s2�V7�-d�Ȁ��2��j�����32<�I������E^���!��HN<�;ې���)ڤ�d�e*3)ָz����1�dQ���00���:��Pewh�B�Y@�r1QP�2�e746&:!KKUt�3�+a(Nt�ǘ�V��a�,
D4�(���r01��5@�]Q���G�`zh�������%vY|0�{�-��r�EE��p�%���0��B?{Aף;O����W3ݪ�j�'tr?��z�5���F<�"t�ϫq"X7�4�
��o���K�.�z{I$�@��k���i�qT�k�d�������.�,�̼2��#]�?��3Y�ך,��I�}�[�3�����ۆ��βm�R2���MH;lu��Ӗ
y,_���8��U@��̀��@�Zu�������H��/�n}n�3Z�{��-G��Ӳ�xJ���Nx�Ë�����R��Pq4�~.'YnQ���넣�Qʽ}-ҟ�i�v�W�{H�#�����S�9e�h�VE�7����!]4��WjUW�]���mc���Ã.w]g�"��|дF�ږ���$"�,M8��S5�/|����s�������,����������_��B��@N���]����RJ�U�m(^�.`���~��߷�/_88 ����=�G�6�:
}�Ԧ_��-��e��I��&$'���5�_��BZ/��H�ۦKG� ��Wp����������� =$ٷ�N'��%���.0]�I�_�NOp�0�S��`X~�2�K/Thhͤ�B)��:����S��3�}1��t��vK���(�R�e�#��_[@m�~Ӯh��\����nE��+��/��Tܻ�?g+F��������N�t:����g��\(��/_h)b\�O�:>�ڡ����V`_�C�3��k?��o��ND���q�;<�ֱ�F��ڞ+�irF��z��ˬ��E�cL~)�y��	\���d@Viy`��p��=<E�b���j�}-<��e�o�/X� ���Z�E�fK�y7�p�j2��@H��
��>�rQ��>R�#��� �J�����`]�d]�U����m�*�+22n0��:�Ak�E��,�t~c����;kp0`�)�ŗ�" �hk�Jd8��2�zZ:e䦡V���Ȱ���0��+߲�<��S��w��P	��� Hem���/?������cY�Ŋ��o
Z����$t�,�,��YF\�m�I�A#�	�F�N��@?��*~�9ְ�Q�ӊ����K�:oi��]e�9��إ�zYFzK?~ժ��P��T����OO��+]ⷋ��F׵! n�rI�����M��M� �B�xjE��?������yp�uj7�blo�~��A�K2��	�̶�fW���cCS����L5�:����D��P�(E��c�:�y Ю�+ a�%>�M7�����>p��oi�ll쮭�#��$�		>���>��uK�Q�k�[�����/Q��7;e��l�V��D(WU�-
3��n��p�ĕ8�/ٿ��{���/6u�yU(�a�G��կ{X���?+��2�=�yT�;%�s�g�������Q�l�h���y��4�2&��u G���O{y����]y|�ͣ[�z`lx�8bi��SvV��ux8uY��#}曚������ͳ(;����ƿc����}yy�d�l�dS*+���n�����@�9��}�:Q�bu4���:���YC����`�(&�cWC��~u�A�����9��_<v��g�*קIV[�n%�򮑢_H�f��ߍ�u�R'2`z�k�M�}�LBU�
p�R���|� i^�(}��|�`θ�8m2�+2@nTF��2V�9%>��f�[u�a���Jm��?~0�'��@�鍩�E�{�_����{�H���-�x�d�ɩ�^��k�r�� �����q2�n�Q���NP�3Q���=���\������u-��
�n�g���O@PS�q\TA"lA����|(]��ӭh2k��Yt�	#G�󁙝�M�7�1y��Փ�w�Ybs��H@X]�8�7��Լ�[,��{6��U<ֻ�ݿ�Iq"�:}�$b��0H�k�;���G������};6�F��n^/���Y���ZY�r�S�wii�&/���ŅYT�)�0�rɓ.ZJ���F� 
(��.�߆�g+����f?�j����jɓ����6�͗�A�[t�
�u4ԿM6��Q�?:z�Ё�"p�0�:�Ѝ?��� O�"2�("Wb�~qd��˖���+D�ȧ;\�/N�8̭��1<�͍�]�-�x7c�z�<���%�L��
�:��$k$_���.Lx�$��| -��u�s�
KH��V������m��WdW����y��\Q��M&a���8J�M�l�E�;P���j['��;���O� R|}Gw�j���1���<ׂ�X�H�+�ǬhU`B�hT7��c7��χ���PH����:.����W���Ī�����869ۉTM��j�[Ȳu��<�V9��5��`�S�.[�n�-�������(@�F:���&=��¶K��tqpɢ3
��)��c����Vu�'�889e���r�>��
��� ���2"A`aQ�8Q�eD� f�k�c`|������e}�r����%�I�0:��A��&0�|�2J���zrk�^<{c���@�P�����
��I�i���[�Ӝ0E�]�x��7�*ol���H���:E4e��0�IG���+A9 ���o���b�����`ۀ;piN��P:/׀�
m���O�?�p.��R#���B��ľ��*�xW)�T E�4Ҫ.�	�]�Ks3%�B�x�M�װ�S��!5a�P�J���Q�p'T2 忬����;M>�'I�_����FSS���j��Ys�/v9 *��S<�?��	K�k�����;�Z��|�q���J:H\�#:��U��d@b� F��ʮ��T�U܂5*?~	͇�sB��;�P�tNq�]�N��n����Pͳ_���D"��`Fj�d� �ƅ�^NA��T <ew<[-^�T���ڹTB^��P�.b
? ?��q_���˃(1�j��S��r�:P�AA����`99��pn�T�[����_>��i7�_��7�ɮ�����[�����x?�`q���'����g͵�p��A|����T� Y�,]^���_����v��?n#�9hP�7y~�����i�Akc���|>
>�1��N��Z�Գ?�0�~:�\�?~���:�rr'�l���!`�s��voTq4��.~�;�npv�e���~���W`ң�C7�\&�2��l�k�_m����|;�R�� ��e���9E�S�P@����xx���Pß?#,�_��\�rܑ. ��A���^.�e8ޟ�yu�v�	���g�Q�lEm�4��o��BL�JN"����(��T7qW;��L��*.֔�/���+m)�(���ON�3����y�-�,�l�~D��* �UW��ҭx�2��ޛ�=�q7(~mT���ƏaC�Նjh����#����=�s���י.`��y�#Α�$�������}�!�v)B<��>Z 166��C&�3�Ō�ny��s���T�`xQ!�%��sO��Gǵ՞ѳ�A��[�]�@���9ܟ�����D�+q�a*�A�yM���%�l�/o,P;�rfJ���
�����B�Թ�u��a�� #X�]���6�-�g��QGy�|���c��J�Ұ�!��Yں�7gm��S�C{{~㨇#*QQ�������c������NDO�'����g�׬��C',�?�n@������^[��$�[��]�����"wi�rN����"j=��~�����nF��^�#w��e�S�Z�9]����}��Ҧܺx)�_6B���=Ju� ࢋ��q�]�B�r)w*�Y\�������5q��-.m���-w�cS�%����Z�x,į��^���LG����(
�s� �!�!d��j�h��&"#WYyӆ���B�v5��36w+�Ɇ��l�˔��K�|Q��6J@�(���/G#�;ǝ��)�e@2:�A����	rb0h�u|��=�WD�Fi����	��}hΤz����:�/q#��bJ�:df��U�t��	��Ŗi�٧LA]~!�2�W�f��}#��w*a���.��>E���L��(`f���.�	@�����V�Ւ��a����s@n����#�`��)-t��v�+yfff�9,5�F#�u�������߹߿.��vgee%�'�DC���´,�I2�8<ԓ�����vφ�5 .�G�Ã�r�s9Kܿv(�B�k��_�
�\>�6hAL���Vi�uǱfhQ�}V�i���P����Z|<��C�� u�H�F���MK��zz�b����]�ȒH�G����`��
],`w�p�r�H�x�ٷH
�{@���ׇ�4��}�|�<��d���\�P*_\��[渀]�w�ýϵ��{(,34u{����r�Ç�(u�ȥ�+X.hOf�cF�n
s��8#c�{������g�SR<��&���X<�`��nf���QۆK�Eѷ�uZA�҅A*�,Aio_	�RA*B�/����1�F���#e�s�%�+��m�
V	�Ԕ�uM����Y"A��x��0�31��5&�K�Ԫ�T��]_T�7�%(`_���5������$��JRZ:���M�S���������ͯLOߚ$U'�� 
�9	(����l���d�;	��~���vV�uJ���`B<;{&fu5����:s��\�O����C���l���E�/?^�+�Ʃ$v�VCok���Hrt�V�6�w \�q,t�Pv'-Y�_�}6�?��"��Kwɨ��8��g�	���аn����V}@�~�S�H� qy��p�kg��˃��`[�J��wyu�M��7�|�\^�r�u��P0��R��H��+�ϝ̥
wc#�k!{s���d��!���_�ږ>� ꥒ�jS�񃆴z�S��4�*���}�h�d�j�3g�J�$�����5?���z��K���.S�I�74A��j���_:��t�*U��g����n�����s0�G�l�����I��LD;��Y�x�M�����_���'�&�/Dr�.L�BL���i���ݒ�Ḧ8���IEI�Y�����[�7+$?��]���
'������m]s�|h�Ii�
@�, xcbx�ŀ}𠠸X�3M�����r������ /S�s��Z:�i(��ԡ�%�z��vz�h�@�n��s��	�rR�8A��@��ܢ�K��tt��#$�d�k*��˯��zBo�� K��'��������ᓱ�͏�>�Ք�?�pzfU�p�j��gF+�{N��5�s���+M�>�"�!|*��-�}���t���Q~�! �}��Ŷ��s��-�������x�����17�K\���ǌ���{c�9���1Tض����
 ����\�ڶ�v ���G��T�a�yaϪ��uɉ֤9ޅ�E7�.h�ŋ��Y�k�^��d�iEmUG-_�a�ܿ 8xi�6	��' r�xH7R@''eB�b� ��!��n�],��_�v	W�ԡE7�����=-�y�'�?DOׯ�x"�B2��V�,T�X�,��ӻƼL/�a�SҐK�y��ʷ�Mj �����	��d�rs�krz�)}��ٙ�Wg5��=^�W�U��
:��)����<M;�l���7���������Ҳ;��A�P��_Kl�?HU���s���`
"*��h�ZD�;�����B���o�y6LN�W0�>��4YZ1�EC�V������μ�T�.�[?���� ���ڠR5 �㮥���E�����^���>�r؍ ��>��ù��*�����v��q��:����RRj�s�1�|p��x����n���saooR;8@��.%`w�W�'�Z�,wҲ9��c���e:D.��m|}g}���Qg#�+!�n"?�q������U#ߍ��0���Sq5����?թ���v�yo�iUU��F�����Ֆ�,�rn��f{3�z\��,�<
�o�b畩'ں��� UlӒ���@~��Q�eo	A]TBr�A'*6UNf>���"m��HT��9xz���ei��~6�sH�Q��..䮮,`�Qm��]G�ބ��g)�e��U��x$Ze��<��"��ٖտ��:^sњ�Jg�_��8��:z�����>��{�z�����Z�-�c�4���+��y����	���,�LH�����ɿ��e���/?�I[��@�HgIҐq�*b%ž� ����nD�T`/���h��"W5�r�% %�NI�8�/��|l������H�x *�2[Iֆ���{3�~^�>����ȸ�#�SG�s�ŷ ,����ڒ�V�_����Z�X�p�7`'gB��TC�����l�������Vuvqc빀�[d3?�w뛚F�� Q6@������@�oj�st�$U�ht�����a�����7�@ܼ�_�8盤�Wיbm:���]i�R���R'��&"�0�gb���E�\BC~Q����H��@����g�����4�����;�����h^z�`tٝ.��+UU��c%Vu���=�>�V6�$� yn�t¶dw����/f��=%Q �����۹�o�zl՘���K(��{!�
���d����c���B���ݵ�;�nA=m,��T{%|3���/��P�j�~�Lv��݌G�}��r�1�x��P\�.��B�0T�L�'XF<�����N��p�j�p�=jѴN���'A�s��iu���n�^�I��r�[�����8�b��Z(0H��ބ��.x>��9j��Gk���E1�Z��بH��#�u��m�����A����.�bUd#1K]��b:���N�ͩ4�T?��=������FH�+ ��ۛ��{�|�Db��g�H!%<oG߭p����ݐ�������v9)M۬����}�^��eil��wVV��9���v�!hr*��,��'�3�8�0Q~��-�x��o����{�yM,�pm��K�J��N�7i-,Ĕ��=s瞧"���˖i���U ���f�S�,l�1��r�P�OF#�[(�GG��U����jsѐ��_<̿NK;շ�mc�p��1ć�bx��`��UFǂ_�'��[����0�����
�-=��_���tSZ	ݓ�ut��|yQ�����1Zn�ST?x,t�/�V?$_�``�8��Y���&�����Qq����
fhq���J��c��O��:~V��G���hR�tX��ة<ՑXċ*� 2B��!莅���! �/L��-,D�����*6��x�~!ۆ��&V�8���m0�F�D�'T�8�J#}>��f�@gX"�*-w���hhC��v��?<T7��Rb����w���J�֭� �bX���A�����b@��b*Wāg� �`)���PV�L������bz8c��۶A�����k�(OJ*5�8㩣7��/=X4�����V\����M��A��U��a� ���S�Ҫ�1��ٜ���_���s>J`x��� �Ȉ��Óv�C7�t����!X���.>/F�����%<����	��������I �� ʰp땄2��"'��ϟa�̔�m���9��B22qYYƏ���\���ڡ�K�eV�jA�<<����#���2;?~0y�=���o������ˍ�(`��a�,��$����D3��������=7���0�FH��R�g��,R�X��2��F�N\[�6�ilϥ���6p�Q(� ���\bR��g�G���8����N�J�_��{�>sf>�x��>�IT[9tt�>Y��Lm��S~�2W�>E˴�x<�$�Ѐ�H�_>�@���a�Cm��M���|6bnP1��_�F�qc��i�4������3���{�P�}	ٷ�$�dߍ5��dI�}��}��3B!��&��i��������������?Ǚ�o	s?��~^�{�{��F9�a�H���u2�n�zuȝ�����U��!r����{���O��/E�mks�7R18��+9fO��wփ�3G�}8�'v�Ν���V��r�ߤ��0-�2��*l�C��DO�������v������y��,��Q !{@�~.��g�yb:#l��~N�����м<��*sL���Je@g�7(#B�d�z�2���m)A����R��$.�P"45?�<i_IA�R� �
��~$"�\艡Ӟ�g���g�8�6b�F+��svv>n`�R(�����x~��fF~`�����6���J��M��55*d=��/�F�D^�����s���J�X���߶>�x������.�P��6.��2���Vю�Aq�#�F��t�����$~�e���,z^a���� �;4���`�̀��E��y3Q���+> ���4��NN&r�������P��.CZvq�ؠ���m��t�f�	W��FQtϸo��.ҭ6��ܙ�(l�.��0Ct	����4_G~�OYOD�)��AL�?(�&���C;}������㬷��ʚ}��{Rg���*��|����%XN莬��s����!~� ��Z��';l��7�5�9���5l��Jx��C�5F�):��J����?�\�����nDP�Y�3o7P$�e&63�HquG��
=���*U�(�.cx����k΢�a��_�$+G/��zR�d鬙�[�5``�M�\�ɕJ�W�����2Sd]�6�r���8b	�ե�8	8I�zJ&�zQX��Ǫ��t.@�Ӯ�\�y�W)V�4��������_V%�kl�R+z�w_Z[;�YM�[)j	N����O�l��q��������u��(t8\��ICE�址�?G��x	� ��l�C���Tc@̭e��}К�Tf$���q2'	ȣ�Ww���,"��2o�^��U3@AxiՇI���bH,�p�ͦ_�Y���N�S��G�����k/*[�P�va�a٨?~Yt�r���QHP��+^�	'�a񣄸e.q� ?����8Ջ|�*1��P����S�κ=�:w� ���h׮1�9?���CF1������0��+Ɛn�*+���M�(0���<���/��X�Kр�U���<��f֥?m��-��)&��� �hI�*or0��2C^4����M���q҅*W�|�!��ƫc��J�'*z)"L��$�dAZ��r�z�x�W�h�kKB{�-����,B8���ip���G� �dέ�v�@�cn^�q����ߍM��T�Ѥ��|��F�H[*�L��ϗ�Ӗ��wrm̅��nI1j��>��{�Ui����iu�<e	<
(����qޛ`�t�3�0"`V�֨�[*ՆH���ۼ����v���?oA���X��K���hdT��s:R�Y�m5��^���Q;�HP�&�e����&����(O�,:���I�����|l����Aލ^	�pF��+�-��|�7S\�hre��'����&>��=�b�a�o|���fl�)��#8�̭ˇ{��KK�7���x,��������c 9������#w�)����\/��0�M��o왛����;����L���S}ڝ bQk�8
�*�V��Sy���&�ه:�%���cs��N�"8�����@�WZ�aϔ=��q������rne��r_���mf��,���JW��٨d�
�����+���r��_�=�]W���p�_��H���E�m�O���͸w����i��͍���5;�Qndj�(�ļ�g���9?�u���d�y��W�B�������[&������H�P)KS�u|,(�E��n��ŝ��Tq#�(���T�Y�g��˖�J�~�Pv�+v���&�28Iڀ�����������1>Q2���I��lF�vg�e�g��/��C���& (]?A�bۯY��(����9<ޠ�V�B�}
�PA�H^c��M?�/�.�}z}ʨa����U�?G!�O��r|[�������J�����x��B0L�>ց��O7��~}Ɗ�=M������*����k�V��I¬eB��L
O�d�g��j����f�&fW�L�0��V��|Iq���]�C2�3<��щ�F���I�?z�_f��=U�����F��Gls?�{ʍ��|�:1�[_��|:��?�&K&���f��$�sa����ki���AU��l�}@̬ll��	!k>�..=���"o{z��x���eX}9�n4����ا��NK���b<^<?�y�!\�Il�|��5Qze�[Nɰ������F�V~��GG+���xI��ˋw��:�_i�7\U��M�d���2����3R��6��:����n��b�Q\���2����<3ޘ=�R=��,n�UO��9�~����% ���

]�G�G4�7$���1+|�ӝO����ϡ�n��?X^]MG�r�s�Tg��^eX��鍻���Dn2�_Xș���� EEDF0O9��vv.;4�>IF�B��wxb�L�� ��  �'����F)hg��,�.mX�z!��I�4N���_*ֻV���L�ĸ4��%�Y�����~�O��{-%>�d7qB �n�n����̔G����yw�rM��Q�H��*��ȝ�*�'Ԓ��{�N������';���߼����ki-|K7SX�9,-���5�qz�f���j��L����ןk|����,��#^��6UcA�U�{p��������8_�bI��x�q����Ĭ'{!E�:BO���h������X�;ifh�T�^P���r-@�`R�0@�����P� 
E��A�:*`W�f݈�����������q14L�~��K�v�mr�����@5k�A���k�L���U�?{��O�\��ӧO�i�:�7�^W�E``*��о��q0��7���5��G^�R4��]~���<M��=�v*���|�.�n$�p[����ёn©5�8�֭[��ƝD����<��<��YYY�r���c�P�uq9Ǟ�_�d R1N�H������CA]�цx����8��gN��/�S0!�OL��N�
֑��#O�����֠Ő�S����ư�z���Iɨk���k><y��/�$u+2g=Z��M\���߶�c���w��)�w%S�u*r�iK�/��]S�u��4���pټ�Qh<[k�l}�����8®;i��2M��~�4rdD��,	\�hN�ʰ
:����C pN`�hI��vt�C�	^W&��hGt]L�Ҽ�~��gda��0��x0����ٸ'Z�S}���^f����z����D�Ѥ���K)>�.(����㮆����
���T����م��c�i@��	d��[�7��~5l������)��-
�01k��'<�Ȉ�i�W�K�Ҋ���O
-Ԕ������XԒ'�n���O G���Rl�g $4,�O�@�_����_�*�#` Ύ�4�#W5���[[%�R���U��
*T�fv�%�_��/w����{��� >Ç1v#��Im7h�[�J���%ǯ����PV��]ҫ��[[[s��cO罂.���5�?1311�m� ��p�� @eKKO�����Z2�(A;�S�ƈ�Z�w��m[�v���NQuړ+�/u`�/�B*�k���8��㓗:��4�'�����-��!/ߤ��(M
����z�㔥�FX�o7�T3��@�_Ph�'s�%�!�om��Dc�@�C��ǫCv���a�{��`p��f-�CI))���M��Xz���p�v�rr�"�K�P7x�����p}/��5�����A|S�",��W�Kn�r5����)�r#��������`f7-q!`'i�LAwx a:k��o��C�i��L��l����z��S�pT_�����0>9��,n�߃V��2��S��3�=�f6by�M�o�ђ��MW��U�B���F����w&7L-,���
й��4{�w����t��YnKQ)q����ܦ��@}�ucB�-4�i�E�z�����CQ�^O�A)��	�ؼ��$5ogIiZ�~���J�*$$�t��U�cwwR����Ζ����ww��p�}����c���12q.�uΣUXT�Ġ]@F$����as�T�F�W�H�)��:	~2�B� �'��i\".�+���ٓ+�n{w#8�o���MO&$�*2�L�W���n>�!�[Vl${B[�<�U�|Z�5BQmH�DYg4���Y5���(�&ի�0}eѼ�m���C�rq�̀NP�%eȁ����In�\𰴱����b�r%zw\)w𽥯/##����իm��m--Q z7��P�FFʠ�������/-1 ����1� �A	��V��3�P}����� q_{�xf|\L�* �@6���ai�y�s@�}�3�W�3�$G�+�=�����9�	v�'>-2��eF�D^�.)?{b�K�R���~Y�U����JMtag'i�zkϲ� � 
I�"��� 	!(��d��N���̔���OL\�7�F/m�m�.}�O�I�FI��3���񀬜����PY��r��-���
iS3t���������������SV)��A�i߿ߖ���I"6�d�D-[9����Q��[�u7i,�������mb AP
ޑ�� A��5��/(p�����U��qe����/{����PFb1���s?á�3��逪?B3�ܚ�q���E�@΀a��� �dSK,ȭ�ͨA�YB�I���N�JI
0�~�.�q���4D����l�.��7��GC�5�构�zɏ.o=�>@����R�	~��s7���_�9�i ��Q�6�Wid�\����нw|R��:ghk�$0��@&=T^Mhj�$1s�f` � %Hv|��WfN�o�:��qc�8P��O*�\*��%<1�zh�-��K/((���摲������O
JJװ��l{���X�����P��M_6���o~V�H����B�9t��N tѹ��R��,^�z��Eo P E���׫�dA �ܞ�j�0��C�S�����q�ěb���2{�A ��L
���>uj��;L�l�n���?ܪ�����N@w%�h{�%l.֔�"���Qc:������TT\��X�U�	���m���<�e�fw%�I������JL�c (��M�@�ʿsA�=����婱�@����(���V�M---�zx����� %�Qkj�6��)����۶��U?��d��ٌ4�yAS7�ɑ◕7g�j��Ah��]����X_w������EՈu*l�%��efC<}�"�����:��w���Ia�DYY�/PlX�����/����*�檝澜\2���|���e._���Ù����@�\�Y*�TV�f��{-GLx��c�/f�_�ǵ�߉A�[[�X[D-�:������	ڧk�[�N.5[����屛�+w��x���[^��Z_ y`@��;6�"�9���P��X�i�����޹�^�Δ[:��ikO?�C�2������3a��U?�*�,�r���܆�Ā�M��ųC,J�T���л����}�����_�R��J�)�G]�N#�'q~��G\�<���ee�j�Q���@فcR*�y?1qh����4;��q���91��S!���Ԙ���j屷dd�US�y�/�d�;4&4�[��� ���=pۮ��d�x,p�X{����OBg'S����+#�������	,VA4��ZV�|��bMq5H6��D)VSKC|��,ѭ�4��u��'{��I��.�%L�֚<ƨCo=��E8�����gD�Jc+'�)�^�6���T�繆B�\(׮��ރW��ȃ�TF�LS��� +�T(�m��q���˓1 ���V1e5Y�x�)���Y�����,	�q�:͑��+)!��%}��<?ur�����Ⱦkn�A,A�7���keee4��������P�4\aec�9�ǣ_uYȎW@���P�ںW�}�����v_�v�$���1o[ZF0�z�Ӭ�GG� -�т�u�ϣ޾>I�X�Aw<���&gc��� ��(����?�(Y�Ir�l�ԟ H	���NQ��bQ�wɑ��٧�|�ɒz�p,7@<Cΐ|�w)�S5�TT�:����/�˃~�z��I9���À����A>WU]��6'&�+�3M>]=������ ,[Z�c���׳��>�
�W�.|�����	��|�DG� �
���nI�;H���Y�
ޱ� �k4����oq�D5������/��lF��7n����y��;�oT{�T�;:"��weUS��ۜ�g����յؤZ�Y�l?�����5D�Ԕ3�z�z44I�Z^�Q.����hdUu3O{���7t�	�Uڳӱ���q�����33����9����Ch�i��[eƜD9Q����V�E߼٢١j��J �m�v!�>�����?}X02S+Y�1���w�)(���=�1�����/.�WQQ���g�$�;h�������ttt 7z?}��A%�	i�c��\�ʾ^b$� $��n�}�10���b����Fbe�}��:�%*] 5@
_��d���oX'�'�~?G�b���֖���G�9����&&`OeN� ������L}�ߏ@�3_Dw��앍�N�´�C�`�>/���s&
'�(��+|�/��~�����>i�J	G�zhJg� @�Fi��ç}^�L�n[���:B�:��4��Όb�I11����z�£�r�vP?���������/z����˗���oyv"��e��H��-�����ݟ��8�U5���W������=E%�l�?xfׯ_oJ,	�FYY[�U30L�' ����ٹT
�Z��k�Yu��9IEwVY>}JVf/���%�ܛ�����Y�����4N66oJ�����nY`hN��'�t�z���<{"Q,�?�R���,�"�,���25͗���E�hej\%��z$���'�G9/5L��J���Z\g���$?/�|"�2�tc��Ia6&L�7B��n��}i����)iz�H!���$��o�K��_��/�p����8�:"�t'J�K-=�?�ɒ	D����{��/Ez��g��-7����9ڟ�f()��蟞fO��qE=N�<��GX;��MM��v���;u��
{�������T���]ts���ѭP��v��\�E�֭���a��l�&�{	ż���
+���&��{D�9�nf�y�k�s�en�,L�E��3�S���s�b��{Xl�,pY��Ҥs��.m��)!A�}�
p�غO\��h�;�M��Õ�� �;��+��Y��L 9��u@t˔P�����ם	�8� &$��>R��s|=|DB���R8���cMMMnVJ����
�����6��n�޽S5�ˉ>6<E��5А�Xd�����������7=�GX�ˎ�U��3�*��²�.�|���
)�;E%$�m<>՗�tuI����G�(�0�b[*�x��,��8ċQ��T�$e��fg�H�p�^�a��a+�74��PIR���2e������g��
Nj�K.	�*֠�t�N����1^�)/ϝ&�h� ���ŻȒ���+��󶈳v�ۊ�r��y��˗z?��Xs4/���Ϸ6\������-�mv����ۤ�laЀ;�\.�п�'^V�TXR2Fg�%A���������,�O�;�
=ۧ�G�w~}TЙ�W�qw,����#B�[8�M��8汱1�ZO.��K�����|����Ǟ��E�@a11���vO�&��Ǳ�����p8��A"SCm���	�H�*�~�S�)�@���ރ��f����D���+N����q���w�`��U�w�N~��f���gY�Wp��>B�B?锉��Gwg��̠�S^��<)��~�hӉ��09H�_�6��uv�N)�����<�<��k2�٨���K�A)dN�k'Y�� u�`oY�����x�_��l��1�H]������Q������|�DP֭��������e�iS�n��574$��<��jo�����e�Y1sXz�W�	S�Mm$5�T4�BЬ��RH7pV;S=6���'{p=��q��(���b�C�u�D�g'��I�Ɨ�i���?����^�K���<�0� �c�u:��& '��T�4��i�����EyʏV�I��<��
��v&y���/mA��w��}� �QH�ڻ�-�'��S�~���\J��}��	�̈�ժ�"�AG �k�K�q����4y��[=}��8��]���(�}m�����]�ٍF�����x����A���_º��$��RЌ��`h�D���� ��O�pI����$^�*��R[x1�7z5=2V��v�O�f��<�8D��������K�dsц'��4��>�u��[�w����쪪{~���J������V�r�!��v*��Q0�P��7�F-�O�%V��L�����~/H6fXի�śW�
&66hrds��ʇ���QP��67'BW�9t��̸�O���V�3��N�4�56�WU��cJ
���o��I���ww�+�	v	
",)�n�ޘ����&��� x��)��?�K����ۺ�ip^������������ʺ'm58�[�]6��k��P.�!`]b���D�z'��b^6��,o Q���A	N�$127�s�Ӣst���F��'=~Z�aX=^�n�/�����[-k�������D�\i�\!��:���&%kS�����&ʲE���R��3�p_��&7�F�������?�:͕�2zvv.�V ��UnII�V�Z�:\~��N���"9)������a�/,���	���{������ҫ�kl4��J������lp#U�$͘��mr�C�лP��A>���6���"�cx��Z�OkclH��{�\�deto��`}kկ-h�C]7���9yvu5=c���=3*`ht�{��� <���QB١1�Hp���'�<7�j�NT�{���M�a��Lh"x7P<<�3���в�X`�"�6�S����U�WQ9#�5�c��8)�aHD�v��3}@�1��
�e�J��ױ�#>��!׳��f-�g�h L��XW�_�s�β��ols����̱�v��q߷o	k;a�/0�hy®k�.G:j\\��o\��>�1$b��uo����3gPU�l��?DyvPv�}o�%S��ۮC�yW�4��Yݛ�ݘ��ȝ��X�����i([|��|�d��e��@,(I�߻�']���/EK�$���� �_0f�Lɔ󵇎8����e��-I�<�m8�"�J����L�ͮEG.z�wWwL�
!�_����ʘ�}����i����_$�HS�
	).����xK7������ʼ��yt8F�7���S&�ir�v���7  ��i0���z��B���W�R��)P��r��'t�̅�x?� ��-�w�V���8�����!V��3r�r�k�@
�'.��0��b���0���DDl��1k>��2e8f�+8Q�Z�w���n� f&��߅�M�(=���(��$"��b���IS֎_T�~Y)`!�UK����O����}�f�Ď���b�2Q��p�	��a��k�ݶ�A�u�OwyL@2���EQ�4��>@?��|�ዏWOJ1��%�ݘ����C8�fi �<���_I,O���Ɉ�?�
���3��|�+�ZΆ�����W�>)����
=^���0<�NT/��k/��9B�΍:��o�C�¨���@���!�Q�Pj]�,����D`0?���2�弲�ȝ\q���q�����@
�lT2@8w��]����ZtWJ�h<HK�⥞POE `$���^�ٴ�NL@�6����F)�֜��8���67�'Ǭ�VJ��[�Db�ЌR�|�<�����ӹ�,����7��F[#z��;���I<����`�������N
���kjn��z"�AM<(2H��9 յ�f�~㓋�e���wZtg�/�ҫ6ܜO��s��[���?��O�VA�I5��B:��򼴽ssz��d�M��8yt����G�#:��b�/��???���V��k�|��;��no��P`J�=uu��n��"dɣ���X���}�+��X�O6�+U_�}�����$$*ob�	sMq����k3B"��1���]��PW�Z�re��h�F�_ �.�C�`����f��?>����+��������)0��w�=g�.|6%a-��m0�v62	���!dʺ�8�Ā�9�zZ�/��*�ck�d2��҅�?|�J�+b�t�ɥ)L~1]�&����V^^�S��_�6KUz�����_/�	�s��l������u>��7:�9�Q�a:��⩁^>h�ԇ�^�d𗾷�"�o{[����/�m�/(���Z i$��݈�g`�a�ꪣ��J`��ǋ/8��YՕ����6�6�P�>��ݧd�Y��i����ĉ�@Uox��5�sz@���Eb(�3(��N�e:��k�5�}|������� w�D�)K��gd��Y�Xc�����NO
��K��|��ȸ-�=z����c	����-�T�f�w,VY({��6bD\��u��֏����%z�ּ4��ڵb����������<�`z`趯��w&�	 x�!���z�py@��Y�9�T4�wz�2�t�ui��\,nG��E��⫍�~G��~���j�)5�̳S�̄��ϸ����f�߂gO���1R�O�b?��'B�䪁�i^�{{A-�+M�%3dӀ�I���=x���}��xeۭ_����a��_�7��$��cd\�$�r�LCe����@\�\sH��e���ݶ���;q�܃t��5�4G�"���P�jC((`�t��^gN����n���T�A��ȟ�m��ίc��y�ɍ�#d���ji��w����=!o;:"�x�3Po[[�u��J�S�@�n���?=��w��I2v�ı�zF�;�0a'Х'����JJ3u�=��M��>��@Մn�d�P6��v�&mƶ��?�����˹[��>E�IV��_l��]�?��o�M5���hB!%����Gy�j�.�[��s�MN�8"�~��;�n��G�>�!�I-nτnu>�ݵ<�� ���|i�]��~G{�}}}�;- ���n�,]-	�۽u�(�:9�	�ek2��e�=�p�v����#`GF����O0�kB�P�ݙӫ�9�;����B,ڧ���+[�k�K_K�T�¯B�Y�0���M�c,ޛ���ZA1k����Tv��#��~��aPe�r�0�u�_ۛz;����5o���}����& �k�����Ǉm?�΍���i1�1WU�=PĖ�RP4�m ׍B/E��N���d�zU) �6�7��J	�O��z��~,$���ݗ�&��r�O��C0w�-�N�~��аKA��ݛ;���=O���s](�l&x�vk-22���S�o!tqf˻f���� �.��Q$��uu68��$��"Z�I8�H�}"�M k7�n�8 �Ȍ����	�A7y?|�4՝�d�H�ts�c���M?a)�T���� ����]0�?�N���C ��D��C#s��h�z��9�����S�q\4z)DN�<������ez�q]�l]�i �*���__$NJI���V�MaB4����ؘ?8�L�x]r����ɚJ��1��Z�gI]c_�8���v�{Fed�R�"���Ԍ�2QW�3f���8�����а�yrF�|����I����yYHy�y�A��+��;�Nn���}q�ps��&	������7J����L�~<�/r�b��U�Qss�Ǯ�T��S҈��:w鐣_�b;"Z�<1Ֆ�+I����J	}�_B�onK�l`މ��H�����ye�*%�>y��h�O�'K�'��]<���iexj>'hvY�n�h�<u�'@дw��K�0^CC��~����>�S�?�/WUU�w��-��{�N��,�� �T�����Љ�����/���d� F�2.�}�qnƞ�܁"�u6��a[ޯszS�d����:����`�x7��z�0
����^Ͳ�9�����@��v#�\HD|�@��vs{;� �	�kqqqv' �&_dd��;��Ufi����n0O��[܏�>~�ذ����d��.M�0J��o2O��d�*����_5J5�[̢�Ǫ� �+M���ݻ�U�u���J��&�>�Xizv��g;vJ�3�8nݪ�b�($D��J�yZG{�T�8�z�y�-��?��QLw�.A�쪲�%�0����4�\�9*U;��b
���"��B�њ�b�A�q��^��Z�G_74��$�jKL��R�71��M
8��B�� ��Y�M��������F=���괅��1��i�dj�뺻S�D�Km��Z�Q�\Q��đ\đ
�Z����\�}�3�`R]|���>�Y���h:v-������F<b�R�n��}���gX6
�~����;HA-|���Tm�?c�qh�R��
������W^������E@�I]Y�˛g��9���UU���_�ih�T+��uT�Z����O��,,��i�A�=d���Ƃ��o��{��j��� yz�}����D�"Wc |0��
��������������w8��������3+/�F�.Բ��zS��s���#J��%#Cf��"����Wm*��y�v���3A�.ǹ8�5���貆�)�X��ܱɰ�rۿ�|HT�Q�M����
��������!���MX�k, ^y�M�/�L�����`l�\����v�E��.{Ab�k>_��/���0����%>�Bݤ��uv������"/�
 �FԀ:y�#G��v'A���"����s?�}���Q��*Wc��u�YN�WK���R����xQQa���d2�ځl&�T&��P�<�k�{9��򧒅#�|���k���Pκ�2L}`p��0��B= (�P����Z������M����*9��-�ƵQ�
>�k����MQf�ܱ����u��d��'i����iw�`��J���b3W����iAa��.cy#�UJ��5�^��P���x�˴�H [��KXBDE�ތ�<�J�$d�ݧKmFj�N e����,�A�('�������_)�<	��!U���w����~nKe$�����Yc X�h%���7iO�U�E�%��-W|��r�.���#�`I�#y����g~�{{Cg��ꥱ)P�}�.B�c׀whh*Ѣ��z�)%��?r�0�ڲ#�'*@����)����0�
��p��E�p�ף�����ax�(��P�1�NA�aU��)̸o�����׺��h}|}[^�:w�����d��[��2�M�:#/�+Sѳ�4�d��=׸���:ć�C�5$����gO�&>R�]E���e=���[��f���8x�a����P�3
=�E��G�ȑ-S�5��hR�7��ӝAQ䫟H"�M�I��7��\�G��z�nPQ�ç�d�i&z�mc/�3>&rK�ӲE����y��X>����)ӄts���D��u�sH�߯-������v�8� �:W���W�.��j�ta�K�oe���0 �  o)'1Y�fFV5_�s�?�y����og5�u������!!=M.���9H���'���l�eݎ��<k���U�3�	3��\�����w�$B�Te��c9N��~|Zsi:!0p����9)����N��x{��2�ǫ�����_��d��! � )B���@���/������3�Q�V�m��q�!a��5QkiM8 3�\_��ˁ���"�LM#x�c��==3���.&��|���(|����]g��r�9�]��Z7�
�S���/�6a�N�Τ��LO���1r��.�\�%�z��L��fl ��wl,F��5]�>3x�M��rWUM
�%y��Sg�W�����d�O��:���	c���E@q�T�in���K��&�~��?~��k (�Om%��sˊ'�^b��u�	��{	,��?IvL�G+���pn�������a:V�����K�<��5��.�X1����Kj�s��]���󚚙�f�+^? #C;ό������?�z���L�����J���2���͒����E~v<*Q) !�	�#�h����utX=�֟p��iuˡ5@ii�G�>>	H$�EZ��Ť�Ěm4K㪓ӛM�5�m��ý=q��}�l����T�������o��v�Bv:��Na�P�:�xŴ�[u�;���3W�EP�_����pJ��~�9��X�Fw"��藍a�Ǭ���&�Ĥ�����%�?'�Tֶ�ce��I��^ON��{�av{[�����'���5�Ӯ�ڒz���	$��h=��M͍p����������2����ne��]�vr�ů�Z�v�~�,��w?����q�*'D�K`�mm�̸�si�YL[��ͽJ���̻#<BN����`	�
?Wpf��D��|P~��N�a"��-��n�V@'��5��[7!��ϳڝ������4���J{f@� �ـ.D���j�&g��n����&VU��,�F�g��ݴ����0.�r�xH"\rm��[m�d�y�a�G�����C-��q���ݑ��7���YXx�.{X�źZ|X�wq��E�#_�n������/�_G�����U�ۀ�~`�(��.��蜎���1Κ��4���x*�T�:]Ġ6������<�,k�kq���$��P�l	q��OB�e�|JnFh儓��k���4{���VJv||\��mk�3@����WV�A�?ceZZ��m�ԎCk���B���W�]O=@Y���t�1>)��uHt�R�_b,z�.�L�C|�r)�����9����gɄz*���8y�x�W;V�P/G@X8y�~��c��rJ�<?������2��n7���d;c�2)�H����@|.�W	��#��\�۾�t�4�D�:ĕ���;m��}�a�b܏�Ird�%SQȘ�1r��(8���Iw)0!�P\�9���e궡�5*��9''#ּi._u��z�y��P6�~HDY��\Dv��3s�_�Y]M�4M��
;�?�P�V���M	F�]�*��g�խ^��1׶��5A�������8Ug���I�ŷM5浳;8�b�|5I��~�?��Sp;�c��_���^j��K�F�Ts<�6|�܌Zd�v^����o��3���:�n�e� ���HЋ��"I_ 9'g"%k`�{p \|.��r�Z:�g8�Vˈ���ρ4�=�Z�Q�/$>>9�b��v�]�	N�02�	H��������,g!�1�� ��\�%�i �T�ù���^M��SS#Ħ��#��\���-9��A�2��5ZM#�cE���/����� �Kb�8�69ф��+�nL���GF٨d�? �*ȇ�XC�|ӏ01�GJ������I����b�<3	Pf�����|�--�ͺ}l����N�-��G��VU�
������F��+&��ԙr뙶����s�*
���3q��Pc,;�NcQ����㖧�5�Hd����M-��k�����Tb�kMo����i�	�i)s=Z��:�]W�ެ�e�C#����k��Ϲ9B������+"��E�Tо7�y規U�ZFOO��A^U��:Uu���(��<N���MR��`����_��¬��?!_�~�lV���n�����1�����؅�X�s����L�?���+�7E��O����?�GN��7g5�X%BSq#Z�����p�o��Hn琋$F���|B�;
i��2��qNG��:x���!v�.�ʤJJ׀.��Q<%ԛ��E�x|�|��N�H�%��Ӧ���%EH��T���Ta11 S�7�Ą�n�X>}z�ڰ�����+���>�3N�uMM��ޜ�Ԧ��(o����l����-�}6�a��';����j	P1Z[[�e��70�b�f3g��v��:9҈Ny����?I2]1@�X����L�?���������9K]�gH��Ot����Ψ!@Fn�x"���A?M�����q�f���'Ͻ��|lcC��x�/�������m����)�ay�Ӄ��6��H��/+ �֫�R�IV!rt�m�"�F�
~Se�	���.Tڽ� yI��om�/8�zn�]E��C�����(o*��;k�9;���@>��G8)��hh��w��[V�]�����Q��HUV"�k��`�U�O������iNU"yZ��Q�Dpr���CVIf>;0h5U�V�~g�i��K�K\�}�[3��]����m��i�-c��Eؓ�LQF��f��oQ;����AJ��Aj�|�߿�xN������"ŉ1)�m4(�[Ԓ3��Cx��8H�����
'q��g-�	���OAV��Ul�pE�ab�5�K�,[�48%���و���H==�N$@!S�,\�M	?�~>^?��n�Euiv��?g`@w��~/:�8�+uU��d�V�4��D>u�	�o^F�LM5�7A!!l�X�~��ۮ��Gk����s���# ��P��bY4�����Smp��g��4yU��]Oy*������(f]�{m5����ed����2-����u�z6*N�:�.��t��p^3�Q�n�^�3����.7VS[��{@vS!�45��W��}��,��)����o7 �9�z	��,,ϖ#�����[ҡ]Q��U��_��f��b\@6���*�F&���⒓���Y�#8��H|�}����������˰��/�zQg�'� �b±�ҕ񂢢P��[�ǌ@�f��w�7'ɇ��~�6x,�T�F�&���n�z��<��	 �+f=��5H}7O���y�R���Yuq���ܖ�ְ[pp�Cc���8K*�'ɩ\�/-��tY�q������7Ƈ�>h��s1�ӈ�l"�(H��R|��{�󳡶k�)�3ѕ��-���_i�bƁu	6�o����Ʈ�o�VlUlnݹݰ�������������T7�$}�KS.�;�q����S`4�˒�C-�ZZ[�zzdѺ�OM���g��3�D/y���������@:`��]�޵�����|�������M�?D���x�>|$�;��r(�������M��7���B��	�Ma��Б�����5I���ֻ�l�-E��[�t�-����Io �G+���?���KM���0����r�bx���Ðh���8�OK���JԿ:������^��D��ΑDx=��%�$� ?9��W�E^^���H��,�U�D\]��I���XZL���l���P����<x��EQ���8���v$�5���c˞��G{�D	�Bs�̌��$��t���Cg-:�'�����$�w�������1��(�@<$,��S�4:�H��O��'v�V�=sB/��p���,�p��L� N��#k>@E�h��j���sH޳�wN��D+�R��	A@P�.���Bж�5���?�a���r�hZZ[�a��mTU�荥��3��V���&q���sgr��~��7��\�K�X#33�cV�E{��]c��U�*�b͚�O._:t���@��������}��f��2{h�ÿ���Xk|��<��z�t�ʁ)O�s��EV6*n��<A����W7O�AQ�-�����gc�܌U.�@������/�"t��"�|M�Hq���	t�����;�����U���{%$I�$3\3#��M���2CٲB!d%d�nH>�n�^)ܐ������;���sΧ�_���1������Q���5�!�ӿDI�k��(�<�u�l%{dR�@�k wv��e�,�y�|�Gmln�9K��#���ё?�9��V�G�.J$�;#�����N �U��	 50�x�93oؿ�Y^S��1����O�9������ݜG�P�z�V�CxK����%؞�-����Ѿ�cI��II���'��� �8}t�r��Aj
����p �g�cZ�A�J���봵�',�%"ۏ2���4:6��4�?h�w���!���U��+��:�*|��o�d�~z�|wbU �};$9�t6n��������O�Ngo��N�����E��M�������&�r��d4Wrӯ;)���n	�R�Q(m�;��ڴ�K{�a瑱<�g~�*+,�>!�u�.|���0�b�`��B��C�m�dzd�`j�<��9�om��w3;�xbbW��]f��T����g�i�J|��)�B�L�@��1���8�'ov�l nq�4�g/85�B��Me_�R?�9.���7�i�fp�Ε}���<�mNW���-2�Q?1��n�)��������w�y�� ]m^^^R3�\��H���0���>��`�}u%���ekP�!�R�Ӗx���|��o�$l?a�� ���m"{?
�ݤ.7`���+W�"/�XqՇr
t@�qS�n���,�7z��2�5���*�3�  M���u�G�z=$��g��vg�Hv���c�a� ��O�<���T"22!����ܾ[( �0��g���֯���D.[��ȷ�W��buea ���a.bktG8��ݽ�A�
�@���1jd��6MmJ��{����hpe���dʒN�C���Ы�b�F:ѫዪ9fyvF�Ȭi�ɷ�	 ��֭���Ȝ�)�??�<������uq�u�����m?�^�����G�W$��~�=�v�UM�*�#--e��v�����~�_,Sc����,K{]�E��nD7
u]����;�I2v��%�eNO����� &x|\8�P�vv����I,rqwl���E*?9�6Y�� 0TS��Ҹ<�&S��I�Ɠ 0r�sH�gyJfv���,�e#����;&��X��eȠ7��agdp~�r,1$,�Z�W�߀!��WU�kϬ��:�I�Sn�؂�4����ME�$��Z�|dZ��rK�~wãQ ��$�yZ��������\TX2�.�X�:/���I �8ھ��G��W&�N�:/.5+���v�oo�H�\zK�^J�y��h~B�ϟ?5q�{��dh���K�o���������aQn!U�4B+���_=�+��U=����9����EHkF�*�ٞr��\��KO��1���_ݏ>�SnS �v��\�0J�R��"E*�o?H**x��������?�E5��S��!�M~�#�$;3���g�����L�6� �������ָ�g�8�ƆG'�?��0̦��k�F�7:��i̡OCBdt����U�SX�����N=9
KWu���P�e��m��P΍��%�w��׌����:�~K�LI����g������x��y&Ck�yt�}�0ir��Se�׺��Uޫ�	b,��w�1{�����nJ��k8��J�}�k�gC�5�﫾S��k����H��p�W�[�(�F�������~�� U���!��۪��J�Փ���x�v�c��s�l������Lul�g ���N֌`+ߌ,�;;w��D=ԽLɕ������j#ɦJ���_���m{%,��޺��8�	|b�j�9��^F�l0b����|�y0��H�V"�-]�N=t�t<�� �^�-]�P��T��,Sߥ�kM���F�ǯQ����=�Γ���D�mZ�R�L�z�J�RZ
��/LDq����}*�ぶh�������9���N��m���/@�T�We����"/������@N(����Ҳ���>��l��y��X=���tɓ�x� �'�))���8� �{�G��4��q���l[�A��)y��̾��A�ZW>�XH���EA�$/���R-��X툚�1�����l��l� ������s�f�0�L2��� "�K�4_G�P�;:׌ � ���T�{z/�����n��_��֮=��i5>`5_�{q���g١�Hp���ל�V�76{�����ɞ$yf^9ՌT*�<k)�ci����ǓZ�9M,���^/9���x7�@`C�fc� )ҙmiiɜ�>f�c�e9Q���؂��/	�gh"�����D5�qZ�&7O�q_Oxl-aS��k���f ����oO/��{s���$����� �<�T��mdnęH����BNv	�
�?�����}�j�N�404l�ￒ<��v߼{�	,��R��*��;���1Tw��B��W5��O����c��,�o��u)n�z�:s�F��^�{cN�ڄ�����u�@�F� �2s�K�LW��d���*�9;XI. �*�1��/�W� �m-�<n��%4���H[˦)^5�r�w�ܚ�����(�fg?�M���!N�1�/���v �>���B^����d}&߽�$������6ֲ�u��:5G��� �n�%e\�+�"P�y��vوt��/\-��*�0�6��Izzy}�wwD4�R�%:��RRR�<}A�F��L�g'�y�c��4��Ȝ-�P��q�<>h�
w^�y�_�;_��]Mu�`�����uk�YRz�4�\V�"�������S!�W�2{T��ru:{zȁƎ�Oĸ��wς P�����_���G֢�����'��gs��Ą���	������y>�Oy�>�lV9�aLxc�SG��u��mEE��~�����(t����#c�|7�{��	� �JC�#�����}ԉn�/�JA��DN�����JI4�W(����c��A�OO����ڱ�L�)�'
�ؔ�g�`���jӧ�T5��x,�PW�aLŲXǊ�m4]��uD�9� p��[�٦������Y�l�ҿ�* 4�A^A�:.51m\���T��O�)�V��YZz���z�-�Nك�}���[4X,6��LJj��S�����扷��6;w���83�I)�Ǔ Z�[Qt.rGc9F �輦�HA�J��n���B���/"d��+!JR5����ࠟEȜ�e���)�ˋ������H����#5�m��LL:eY΄�A�zIf��&��2~���������k��*S����CBv�����6�o���A�N���N$ob�Ջ�����������j�'�����s���<d��X��s7���S0�E_2L��^�}��GF����w���u��^�xWT8Hh�L�+�ã�����F�~��D�r\�o�6�t�b�D��٢'�����w+(��|�^�G��~�X$��a{|�G��*ێ�ﶴ[���p�<W�2�D8zE���� ]�a���婀�`��b�>
���*�V�Y\������\�o�r�����x��w����NMq{=g}���#%>ʧGBAAQ{#�V���s�t���ŋ_7L��i;W0��?{n��|䴜(�������2]{{/c�x�*��s���C�/Gy�A����%�Jj��3f�ra�ü3�Cn���V�sTT�Ѩ���4K#�q����l�P��e�e���1��s�F���U��9F��ϻ�xn�\��|@-$�vB5~����}x C�a����b�,,��e��m�KR�(�*���646~X\�!�m�c�䔽l�5gZjc�㫏}�r߻Շ����y��x�O�"�Q��H�'�]�ep�x`�k
9��������������U���y<�4��Ī�1��Ҧ�,�I7&�J ���}+��s�ė���Ռ��4�[�� �v�[���d��9i�̹&ɋ�|��TȻ�s�K���b���R*X���265%��?Kw��ʊ6G m����o烠kD����y7��y�#R�is�o`v�ɼ?�a�a��a�<�I|��L����8��r��)@f �j�'4�%���+�����o@?D5#ǲz�Roƕ.JI�ț̬x������<S�`��D�w���5.�9�z9ǜ.�l���r�8RIpf�B�������������N�����	�~��͸��ѿ��UUc�>_c+�ȴ���;�-
5}���EϷ�4o�WWF��>���<�H�[���uO�I��n8К��h��SBʿh��o�9�v�5h��?>M��/���?�\<�p���/�k���m����d}5C������k�^s!F�$����0+�T�'�}.]�|�E�~q�g�̟���h:�@ٰ�*���5_�(cQ�f���d!Q��8MM+����C��^��E�q��&���5fw�\n	һz{�*�Y9yx�]k}�������zڅ��ׁ�Y�����+%��9q���A:g��e���e��Z�W�a��b隠��E�W~�YK"=A�_� �s)���e���nRbG �[8��)4�]�9 �x׏��F�TR�ޓ�^��QCJ��T_$/��6²			�{x�#m�d�\Q���������U���/�C���]H;�ݩ�##S��*��-�B��>8_߆�=��66���ؼ�j�yyr�K=��ov���9^��9Q��=�_��i����ν)�Du*U��"� CT�U�2E��J(���E��2�ْ9���=�-s�N��b{j��i��H�B�
nn����+f�sK����4װ����#�����-�QQ�߽���e[�ջ���S�k.�����T�enl�tv��Q�� ��:��-��8`~���͜�������y7�������%���A��6��*�=+e�W�0�6�Ry���e��>�>=�8����0��kb���[�QiЖ�Z��6*EF���}����C���PG�;nnoj�&=
V=S.��1�z�Ї��{�ccn��Ky�"��eqӝ��?c���� ��=�8�B�[���i�zԽ�݌vـ�G8\����g/��H��殦�Ȣ�x�.G)��˽��֚���yԁVA�r��el�6K@M]�DĮ��[�8�u���9�Z�����]M�]�2fBY	���Kӕ��nm�9�ėX}�}�:��af3���U���8�2���j�VH;D�zg�1$�I���A���ʥ�OF/��ܢQҡ�@#����i��(�4�M�9^�4H/��Q7[�X]$�!U�n��gLĢ$n��ܹ&ԝ� ��t�jgz�[��ϟ�yIxU�\w���my���^ǶࠐPwnR��[O���_��PPs�̝s��������9�i1"%1g ��P��m*8�#�a���gyKԇ?�:^��;Ҳ�(�i-�(�pK��z�� ��Ksi̓���C�F>aR�����|�P+�O|ӯ��1 y.����j4�hT*.���{B�# $�><��C7;��~�B6��=<2H$wN�>��#�?���J��5:4��G�E
��C��E�� ��I�����4�R)))EI�{��d����\$D�h���������=��=�ǫ��x|sBj1%��ZhmP�"L�G�)��N��./<$��]{��t��C֡T_�>�B���K��Zt��������YH���:�"=犟5�Nh�Z(�����@�{{G�oߦ�@s�Qf���r	��9�
h�z5C����3 )e󍅭��(���σ����c��4�5���k;��X,�V�M�>EH��m��͹n�&D�����G���q��7�ϥP@��AyO��H�h�9֌l-5�)ր`��}���7�;8��2u��RV٩��KbL�=�)!-=9q�\�����p�~�4����e�|(M�k� �e�\,1�>>���Q,����$3B-��}TY��_\��A���ҕ+�[��-w�غ���H k����6J�4����7#*#ceGM�_o_��kv�Q��5NR�R��=�\��a!UK v�����Q6���� S.����{�I�	;qV�*�����*OD7�SB٣�A�M��M�����V��#��7��s�\�_��p�^5d��X�\�Ƹ66$�)���Q��h���ZB�z���z$���A���QFbSW[��d��IͻZ��ݵ5aaaP8�G��_���S���$�����[?9&B�>�o��=����<==���Qዽ�e�]{�t����������:t��L�u�q���#:�����1'��G��>�}�B�j�n�	��� �=�3R����a ������υ�U�n͹K:��d�y6|�u�h-J��R���xb�sm�,��KW|��%�}�*0p�Y��e����@�r��0J����c��}�s�gg���~/�olz���
{�T1t�E�[+g���C_��L�v�V����w/+�˥�h_��������4J��5��*��������w�ZB�<f��;���X��!mTH�>�^�k.���(��������7�7-w�@5��ǿ���#>Rn@���@�H(gB&��"OV��4@�ic������.;i~AW��º$f�>���A.߾�b�����Z�k����NH�G/�H֌�,.���ArK��ؘ|e����> Q�f���>s�o�(j�C�TyW��s�Ld�:a1�S6���R z��￮m�������^H5�%��B����
z���c-��-'�r7;��G�o�Uv��	7�����*�ں:7�lĿᗝ�*l/�-���)�᝴ް	��˷�2��>�zP�|�� �l�	@y�X��}�Gi��KK���"TU��!m�ޥ�p��4ܡ��m�d�{�Id�����Ş1-�!R��~����$9�}-|�:@���a��c�aM!�s�^*]�Wn��Z�R)�����#@O�L��a)�Ť�qx�_�,Ss�Q�zʅx~��`F�؛�n��=U�?���<��E����o�\����y&��Ũ*�
?.���N���������+Fy*���c�y/�Ȧ��Yq�[[�E��Ѫ�÷����U�I��u��P� ����s����ES�����9U�'�M:��.����٤4�zђ��u[+��G��v��� ���fz�Z ���T��@yK_Ň�4YQ�F���]Z�=Bf���~-��op}x�<ћ)SӘ�rp�A$~��x"T?|��43cFP�W)���X��da���7er33��"dܾ[~�ڽ`�>-����f?R6����L�ES?���ݾP�c�oO�����c�㬻$R�5��ܳ!&$DF�;���B���泞��mmr|��bY�AWFK�*(f
�>��=�ҟ��.,��i�Z��)�A<�\�$�$�+A��~�G�(�DA�4�:�J"��k';�@�0��R��TFF7���$���]�"<GW=��;���2�F%^k�M�̻�#|s�<2�$���oi
y*���'��h�H��yb`4C6����b�H�Nii��@n��ܿfQ���}x�A��F��{Ș���T�}�3'KJJ��~! �M�����]<7�B!ޫh"x�� 
aD\\]����r:�y�������<T��=�n���	�S=�Κ�G&��p9��U�u�#���7�brk�*U�#�%���~���X�������X�[�5���|�ds��n��p���t�xr�?,zZ�۳tYۛ'^�ʠ�:/elf�;�D��R�Xy��aN�&&ӿӦ�r�=c|�gq֍��W��'�z�
�o`��D�x���(��GB��J���8��oR�OI��!�82�2��!�k7<����9ɩ'�	]����Ty��z@}�$}^s��k�y��컦��W9��7 ֢v��=  ��[��J:ߩ4�EɎ�(��ۄ ��]	Cs�R*R�Nf5���0����sp�Ё� +{�-�Ħ:s�θchHVe t[�%�[��}J?}DL� 	Fy�-F��4�$RL-��>*�ы��1q���jtRAq#@����ne	���z�,�Y�BiJU�C���p�����1�v�� ����O�Ɛ��~v�f�L���eh������y����s6�ڟ*3�`h﷥Sg��t=U"�*f�.X|���oF5��h��=+1n�s��*_bx�L�C��"�$�Cx�\�b$8i",�	"sd��l''�9c��ûl�!N\��~Gq������8IZ��~�=�m���%�Ɏ�v��=�VW���W��vV��lXqqw�X��W��>|�G19Y(�]J��ec�r"��KH�W��b�P4{��y�Ч��Q.��T��3
E�,i=��'�� � k�E�(�򬌅�<��lA�*º����)�����Q^��Ł�f��e]YFrĞ�|�)��n�43����#3�����uY���%�Y�
&''��peh�L��F�r��ǐ�Ώ���,.CD\".)s��4�3�U�xe������3��	���'!wh-��Z�+�e�h�.�$�\
�@�īv�&��)axg�4��T����O���q}��q�g{/������3e��>��^;;�tE�̛7®�'C-��1ǋ�$�b/æK�v�hѓH��<� ��:�$s�*E�������'��^F�?�a��:l�ӊ���v��z�#�s��q��R�����ݷ�Rl2�����{�	kB��Pc+�|�T�0DɃ�^	Vlo�������b����7��P�'����k�E;�O��{r�o��4G�Z^PS�ݩ�w��o��:O��5Uoj.544�\���I��l���n��HV?��ə3���"�CG�!"&6v{5��^��M)ᶏ�:h	6y�T�C��͆��B��~{�߮����>��k~s�9����ȧI��5��hWuu�X��߿g�G�[�]Y�.t����M�Q��1r�q/���ĺ���׳F��L,zZh � ����9�a@kԉ�y�睏n�v�EEӻˁ!6�v�Dw��!����,^��_�
"O���:�X�]T$!#3%>�҇���)�cP��.�8D����Fˬ�r� �%ؔ�3�!ӓ��R���Gꅖ�Z�<�<���C��4�R���w�������M���\�m���B�^M��r�q��jN�@�����ͷK|à%��7d"�SX���	�?�`��3r��ǖ6��� c��-1-�	,q�>$�2���;�H� �}U�\>5��P,���pF3f~���	���pUk�� �r�x��p�U�u���G׸yKyK	����?Vy����T#�����8�3���i�9W�T;Kvzgg����$���hŷ�q��?Kcw��.��V��͜�E��.6ʷh�!:��`��M*b̔�P��"��2ҩ��pv���a򡜞^` R����������'�w�^�9O��i8x�7w�T��9��{�/=Z睟Fq���>n�����2���=;���ަ��C��g������L�W��|��������(�&?����ɮۓ��T��4���%��n���8��-����E�Va���?�{b,<R��<�]������&T��� il�Hz����[;:�rtVO/7��?D��L�λ��_�[�5�����sx�>O�P;%��n�����v�(O<)�wN��Y�D�|��T�'
�,T��\�G��&)5]>��A�g4+�%N��S�A�٢]�)�'8���Z�΁������wD9cNV�~] � ﲽQB��qj��y+(����	�:�C����}�� i�gC�K+k.�Zh�I.C�V �o���H#e������888��{��E��/zά㮸H��>J��95uĭ��J6���f"���O�������)�S��-:�B��������lP���q�Jf�Sǵ<�y�����O�Vb��z�Id�b�h�A���|
l�>�MX#ˉl���U�(-�xd��/�=��7�.�Ą"ύ����A4H4s����hí�Hv�j%��7�t�������O��{���5�z����` uδ]��;���;0_���&�g�z-����%~�Y��q%����TĖ�ϻ�f��>y��٠�/���z��}ґ��V;�����r̵�����������Q@@�C�"�y��BUTē���_g̱5CK"i`�44tϟ}о��ۻubL�c�pZ��aO�q�B�E��/o"ۓ��Q�9q�Χ!�V�N꘿!��ʊN/�<
#bI���LN�) t3�.���8��Ku@6�5�#C�u"�=}�/��!Js���S��{@z��y�A�K��a���i⯬�!��H5`5dB�zV	��,�_��	2���</���ےC�=��Dx\���c�9+����˾&��m]]�����ѯx-.v�"^���u��f6
~�N$2~6H���~0I���Z���yņ�?�H-,I}�IIdΞ��Ӧ�bO����<�_�/���� �x�ÙF��V6��I��Gয়:\��G�i����tTU�Q�Sj�.OMj~�Pe$!)�j�VBi#�\��vQ,���\��tsg�fcD���)���>�6�`y	�{��h�LT�[]��Őc�f3*>��δ�(�w=��^J��	�u�މ&�X_����s��ǃe-��ς�cd���TB�l-*>�Դljm�ս.Rv�H0�~�y���!w�X��sN׿iaF�d��
%On�N�x�\e����L��|�KW`�*S�a�l�B�г8���Sǿ��c��5�V�IR/�H=O��3t�Q<�������\Xa�������S�-n��\��B�K��IP��m� �&Щ��n�Ik��*�����fV�J\}�����/ڋ~�+@�7��Z���YO��便�����c��<vuuM,$`�1r���T��O7����q�$]S.�NN/�2s���7dd�A|ԀmwƟ��9�zI
8kA���B \j4���e�y|Ȍ���Zc����+a	�\��}>���~�T�������i�D,1��\4'�B/���}�{�����Y-/���u�H��0�Ú/�n�ꨈ�+Av�T^}���BQ����v7���y�����W[i�RI^�Y�:= 򷕫O�i?�G�5�nʠbxi4� �HIz˿���A^�#/+<L��M,tl'<�4���7�Í�!T�1��'??�MTÆ&�����P������b��CflU}�Վȷ쾡G�}��_�`6��Ў)�m�L��dP�l0�땫�����Ӧ9��`"�;�"�֢O��k
+��j0$�<O"��!��S�޾�s�ϖ̴����7}1�����?��NI�7�<&{��W�Ξ���>���d�tl��\�ׅ.\��?��r��Q�ԉ� uP�~vF���fcN���h�j@ �ܧ���0����؉c��n�~�7@��MJ=��t�9opm:'�yXn��SݹS��z��YGW��:���g\y��;�R����	�D\Kq1.��s�$I���S典jl�����%��0� ���n��R��k�w��m�`U�`s�3�	��~�3��ٯ�x���G/���&����vv�/��z�n�0~���m͈��RH���Ej`h�;���,"����R�.y�;�������5�Ҷ6��C	�4Jհ�{�����$(xk�GH*\�l����ec��W�b�����FZ�Jj���ʚYX8E��>�z��x�-2h&^�8Gb4FP��
����.շ�HQ��l�>���"��x�-��a���?G��k!a��*=,�oo�HM�Eu噒��^s��1w�����Inv�}J��꾪:$Y#_�i��|=r`�.�F���!�h�7.9��1�"�߬
�Q�P"�ҡ�_�UF������XGU��W�����uf�/f��?��[^�PzM�H!��އ�O[��Q�go��x�Q��2�T��t��鯤[,�r�$�>,"7���i�,ˁ��(oﯸ�_`�C^�s��WINՌ����#::4a��P���������rW��k�k=%W�qd�����\����WMmC�"r�����:�v����^���2�Ts����GAlQE�k���y�V���3�I���B���3kkt~�Y|�γ�z�1S�Oo��sʾ Zg�C��*��d��������-���M�E�*M���
�_(i�1�W�eukF���}���UK_��y�x�t�)=ނ	9�����e�0�����s#5oب4rl�]�F��p��eo�Y�]�v�%t{��j]�������l`Z.�o���-��7YW�)u�L���\������f������(hPd���Eů�P�8��Z�k��A+�ޞ�[X6s��xK`�Vvt�u�[iX=���;�]��0�u�p�Je�5�R�`�b����oC�cD=6���y��2���;���=��P�u�,7EY��~��x�����U>�o���/�5W�#�7*�k���������U	�awo�T�q�=D�+��7Ǘ�s���=y�|h�ݳ�-ON��)+-��̌�+��;��=bb.t'��ݖ��ܼZ�zQah��E�W�TJк2������Ӡ�@��K��T���ہ����:�={
�Y��17E,�xb��0U��lxg;Ǣ�Gs��QXC�3�{5Q�9�G*+{�H�M����ÖG�G�(���p���
"}�;�ǅ{{�tŞ���c�
����>��9�O����>�^K�+�����E�����nHL�`x@�&ҽ�`mxТ�����K���-�t~˔z��ݨ�w��3�W��]>��y;nu���e^:w����ΉrEZ�u��K�<�9�>	P[��ޛ����|�'ǈ�(��lq�q�2�����O� %>*'V����r�E?��Zv�
A�񴂲OȨ���u�]�7��S��햮�]��]Ѱ9�!D)�y�i#uL�4�C����|o��	�����p��W��ǎ݇G6�Gf��<4�U=�r�)��+&"��O����4;�l�H�D���BĴ���ciW�i���׉
�x����������g�w��ߟ|���E8�y�*��e��b��mQ|���nT�2u�/N-�8��DV/e��AV'���"�\}(He?�0?��U/��h��{{{!���*�_�h��~��? �X�s�����4���!W�����K,��o���dc4����]�o�s��l����mFDs��+����{�p����e�
�������FZ�x�>Ř��V��$Z���0I���Hѕtr��o�-D캦�<O� Wf,<{�l�:���KQ�2����kT:�ݳ�yx;��q���<���v��5�ޗ���=6C9�C��"o�p�Ցa����i/�}��Ἳ��NfO��P�`Zj�@��S��� l��3ٓ�|�i)t�������� Dy$�����|�)������2��	.mB��u���ۙ)t�#=����O�<F��S�64�Vz�+�/]�r�P���pJA���&Z7��G�x\����H��2~��IX�&��Gם�TѧhTI����KR�F$�n{�ܫ��&8h���j��I��H�C҈��a�P����bKs���~���F?ۑ^5���*V��uI�+r���2�K�����n�R���w5}1�O���˛g�a���/o�4z��5H9o�>~=�&���,��Px��� o��2�E�Q��G�nRo�qxyyk�X��p��EZ\�wɊg4�OM�/̎:]�����Jn+މ:��������w�Iꖁ�e�
�_�4�^o�X��n�
����`m����(��2�H&�p/얻��ȺϾܼ'0R W��x�/eV���&������?�f=��۷��aD�VUE(L5������U%�]�+8=9IDI�D<�̂vE	՟3T��)Ar�W�1x�M:z��k��M���1=n��ѱ���|P7+W��ip�����o�Uo~r/�ū"ss���i������w����_�V��m8�-,Ш��L����뚠���'&��+���yΫ��@mz�z���Ąb��ڛ����{�{�����|s�5L^~L�� NZ�f�a��]i�^J�I6NN.��nd(������|d���:� @��o��ze�+��
@Q�������:��!A�����/\�;�M#��I )Ҍ�)E��7�cE��+;��Q'�F��_�9"�m�����J� _D����u�N�E���*?j�����;�W���qJL���♖���ݠ�Τʨ�9`�����tQT������~=l���)�+^0(�&�g�:������̏��e�Q�i��c ��Ҙ�G��� 5�mn9��FY99Qx�~������:��ӛx���xc�֖�Q�Y�B�?��#KKO����)���u���m(�#�R��}/}	ZEW0`yZj��īu�3��6��ܱ�u{?��!5|;�n6x�����vM�v��5������=ы�?.rTs�$�W�c_Ot����)��il���T���]]�^ƾ��"�;�w� ���nD����ؕ�Ţ�kj�aD2K��e�p�U��i;��:���gM���Ź$-��$�Jku�⩺^��3�$1��Bl�?��z���d*$$��^��(���hۢX�*� 6�;g@���s�u-�_�V�2R�Rg|��W����߳MB��I��I��S��ȝ;��)�ߊ�v�L�)@w���E1�wm�I�b¸��͚fW+�t���
Q�Ǐ����)���O$�4��#9�3d���Kg�#z��
{5����G����DPQ�Sh�0�	#��ߵʄ����%�j�D� ���2����s�N�~�`0����$}�.]���U��z���t�[�9m�\$��p�����L,�?UԿ���X�ۂz�;_{U�
�GR��`�k�.{���]q[�!૷���}ۋI��J�N�Y�S!d��v*111��@�%�w��}ԥK���w��R��� f���W�kk�HP[�{��rpU~�����D�����'we�;�z�4�N��F ��g��$�D�@�-�ȁF�*���+�6"W��s�ĄM@t{n\�_|N[�+/.����Dn��H�%��Fw������m�?�ϑ
!n �z_���fN����e|�E��&��#��X�(ص
h�aV����Ǧ\��rb8����8���ъ����0OS���&��!����ܡ���`҇�j/J�؆��>7+I�:�����ss�Oό$ugSFK[���u<H�M����Ύ9-�CJ}�m,Q�,ӡ=��u�+�%D��p��(�_��k�T#w�c��?�b�� �i�3֯������c���y��꾖�>/+��o!������S;;�

�E4�\�|�"s��<�c���%�ʅ��J�����:�/����L?WOb2�m�3ر�x���~�mK'�B.�W�������r^[���o�����D���XkÎ�i��ץ;>MOKKc��3-��Q�m�ec���k�����y�k��F7ve��A5Ci�&X%�k-u��H��.iEE���N6�8�UK@��ܰ}m�{$��I~��󼻅��1ᔦ�N��G���Z
�8�<N���P1���/�Z[#.��	��TXݞ\ߙ\��>�V�ks��)����Wo`���J���Dk[ݿs�_^��u��l;I�fH�~u�~����P��}�]���.J���g�J��� ϞR}���'��\a��)�-�<��Oy]��/F|�ȝu�JH����/���tt}79@���Ni��`(;A�;�����V���|����"�O�i?[&�raF�@L$�W��!����h�-�?b_=�q�exD��ۂ���(�F��]�M�[�IE%+M�ڙ��3ݢx���X���\<�y��<�FĂ����W���y�Ju4��}E�_�9��i�c�ַ}�"��%�,�H���ʝ��e�̹�|�c��^�Z���Ž�IT�\;2E����w�D��ӳ��"�X����!
�	W����T�B�`@0�~J�YG� t���Q{~
'.�&Ǚ��r��w]]]��7�s����_"]�z	/zץ�$[0V��9؉�L��n�~��ѣwp���]Ԭ.�}��=�]T �$$>�\������*�|>�#��`�x���)��ڱ��ص��BLV�����d]i������Ab��臃��XIM� ��h������3֞�gdM/]�ߗ���С4�vF6������q\V��mU{�'��������I�'��t��3�7�cPZ؉0��N�c��#e�&Dp\]/h����� ��5��:�g~^�%�m�N���'��R cᑟ���m\��A��,����+��Ñ[$��CDi,�ߥ9���x7<�	�`z�+(����_��,ͧY�t��������w��.Pdɲ�lr�NM�$��pwo0��u��{��A�&���Ib�-��AY�-�	�p���v�~�f���Jm|���xE�C�3����g@t'#H����Av�8�At�.�7u����<Q����^T#t�Xms���0��u����u���v����*nv�&:%�raEZ���XX"��=�42��8z]A�rԳ��^��Z�gh�[|�.p��_��֍̒���y��#�!�����.o{�n����S�Jr�1�<8hFl-0'ӻ+%!&�}��e�g���:�$ȩ��ܾbm8Ψ�j�h��r�EE#����=��"���,"&v�� ���O��{=A�R�ib?��_�H��YA�����{�1v;o�G�Ȇ���I��e������f�{y��;�op�f���2���� �B6�^�s�~ّ��7��<e�����)-�	9���W�V�TBT�p�2���M��%�����nu�x��}@hη���>�����rn�}C�2xl�(���P���?t�r���pM�I��a0�	�)�w~���ș�r*��I	�+�RS.��G�%�Ƚ��c����_�x`�X��;��4䮫<mW<�5�[|�h��F:Eѝ������/j��
[��O,w��H	��*%vv��6j�s�S{uC؆�Y�<S�ck��f�y�~�5|���Φ�<��^�3S��>xŮ\�-/���+�Qr6��/\���a����`8vM6�siI�@�k�M:����&�鰥�%?�p������8�[qY��r[�Vg��x��'�U��ʫ����m�;�-6-� OZ9��:D!�
\o�ȢӶF���3�;/��g�J��Cdx^�8J���"WzO�UfP�m^C����[[��(�5����s�d"��G5� %��(��R|���ff�k ��j���<�H�u�xOvw��a4�X(�GT��_@ɛ7C�ẂIo�֩��J{�^g=l2Ev}�Rz��t��)~~T�P���t��]̌	߉�U��"O�W�l�;(�|��WO/(�u5�s���s2�P�V2�7e1�X��1�{�+��%<2��!]<7.���fy�	&���QdG�h����˛�"�����s�\�	�����;`j�N*0�ȃ׸t�^�ڎG�1#�/�=�+�cs!(rS���3����yDY��ڬ�"8&������S�j�Ґ<�;<Lb,�R�cTYZ
D�⇶6+3s���wl�pT�ֳw���q,��IVK V��.�ۻ���18;�?\j-���m�dvfIɩ��$ǈ��rs}HYF(8R��1(w�'*1!b�NW�����<��-!���}�(�FӋ��!����"B�g�H6��1����=�0(�XN9��9GxԐ���nU�Rd�ϩ���J���(,��b	]�CFA�)���� �m�����!"|�J���I?�A��0�	�H4o��-=r��Ŀ5GF���!F&
�"�範w�x�P����Ҿ��\�|>�Pط_�fz�7��5ց��[����%N{�'�u��}�x՘�c�z�S�]0�{��G�TBQ����ɭ>d��t�1̾Ѻ�a��)�@YTdi5�Tڵ��~|"��0ӶL"k��Tǵں:e�$?����O ,����zx,����RBe'�HI��PJv�ΖU��3��
!{e\��I2.�2B�&�����|����qw��q����|�q�gˁ�\s���3ˮ"��ñ�/�w\�WN=4�[�w���R<��'�Ali�-q��4L����3����|6����w@TN���9?��� ܌����y0>dN�����F��&���FZR�j��j�`YV�f��;��F�N#K���f͆ƞ�ж���r|��m��^��_��2X��C��/,�X��z.���=q�k���^��� �voHepӷ��3�x�ȃ�PLg ��Q,�P���Ґ�vp�L,IbO��~qdL,�KS��&�J��}��e�A٣:LE^���9�M Q_����m��
5�?x��="�#d��BYp=�+Z�`4���PUZ���v�A4���!�Ǉ��>��cR�jV�{2ȫz���?�T�K�d󹗭2w��i�m.���z>{���K�P#�=4o���c��?~-`��y▴x��%-���������U�pk׺QP���b\�4�4�̓�At��nq�$�>�͕�f �i��&�`j������!b|@��N��F h!�$�.U^^�`���[C���!k8�l���%'�O��[�΋a�m���m���Ӿ"oem����76���W�F#x�F\=_�����w����t���;w�u&��/���v�K�w[T��e31E���E���j�|.*J���-J_�y��I��T�)5������EZUu�O-id[_�j)�U�3�N|}|�l�o����qV�:55uNSK��er+s
��j:5^w����ъ�H(�;����� ���Z�K���|�P-0=��HNª�ȍu�z���5��G˩Y�þ�ö���>�y��A�UY�����J,L��!R���E�ww)���l�������MK%u�F�!򞨻i�����JDee����ʜ��`�N{[1H�'���������n�5��[��0�ڃ4��Kn���=y�����6��>�	!!�@u�����i�����t/�3o�s�}�8Y��<{�J(�%��Ը�*7Z��[]9���\��~	D199�S��	Q�y���R��v!S��U*�9�
�ZR|�'Z�WV��T5�3Bڅ�b(�op�BCK+��r�P�ZUٝ�D"QRZ���W܈JW�1��rN�QdM�!��pCs�-�"�����$���dX��"TZ����B����������K-��e�@��2U�8�REȗ�j���q�w��ՠx�&�@�Խ���%��W>��^���.��q�W"�����S-ky))uuyEEC//�荏��ے��<uby��+�HZ� ���8�|�SP�0��~94T��f��=�<O��{�m����	Uh��J�G�Q2��)(��3Y�er~%�ć̜�;��"�Y���:F�~��[.N�W~���r�nٶ$d����pF������Y~&|����|>>�s7�̧�q�*.��$	�K0특gm���u9���?M;d(�6�u
0_C��eSE����}6�o7얦L�
�x��iS��
��@SWiJ�����\v��^��sp<�N���U���j�?�P~��ia��+O��-��25�����&�yq�U��\&�B	S<m��^����[6�B(MN*m���]8����F�tӃ�����K2�$��������c�g�$^��*�ѧ� �xmz���̪)���sN����ww�L��]��DDD�5�\WTf�F����cU��p);��$�p@p�����N�y��h!a��ؘ�	��VWC��h�=���h /��.p���1��:���
��^��ӎ�vT����4�?ͥK6ږ4w}�AF(9ٞ#���'���������k<"���J��쑗�ކ��a�ݙ�;�� ������S���l�va����s���_��U�kb��˵M���|��t�+'v=̵-���8�M�\�)���I;'�o��>-�a�J{eZ�����)i�2'��}d%���}����I��Hq�X�ֳw@w�.M��$s�t��Ȋ����QQ��$'add�g&'���O�Mk�f�T���{YR�W�5wF�-@���TqqqāV�7T+�I�_o�y G봺#������$��'�sJ�T��a�F��-P�w#GG|4��>)�Is��^�11~�����1ί2�)\���ʊ�Ҥ��?���V6n:��(7���<dg/�{���'o�%��5�!��Tʻ|Zr�6��앹>�� .	��+���L�}��z���7X<l��8�%%B ]V������~%�lX��C����Ńmg7~�,���kHE_�xꜝ:p�}_�uO�C���$��_"{5��	1����ȷ|o�^ ����"����T����Ez		��R��|�����^��an�]:)�H���l�3r�we�{m�����Q�VB����nq��A��m*���|/{zh�;��j���C4���'^^'pUL*f��nz�9F����Ĭ3ŝЖɦ�=����555� r&%��.�J{��+�Tc3t\�*�ML�,jci��,�c�{�3�\�o��ɮ�q}�fWÌ�����g�e$㘽F�=���va �w+�����ݼ���l�Z�т��?�W'�[��8�WT1�!�Ȱ����`��d�9����nk�׊���C{���OC��`���L��ߐϒI1ʂ���Rk풙�N����v��z�e��zz4�y�苈����~W++�Ț�Kڲ<�	�]��Y$���5
.ęV���*8�3�߱lu�k&?-idH�'Z�ᄺ�5�����;����ыp�"΂��}vj�7�ODw����~���iE�lZ^I�	���3)K��ic'�5mkI.��ܶ=�)�=�g"���v}=���я>�vN��K߀͵4����B#L*,=�B��R&��R���ǋ�~���Y�_��,���[W�h�u^��Cd����0�QX	P�.Jq�?��F�%����t\�����������L`�]f-��T��l4Eh+���)��cS��Nlmo���|	i�P0���܌���Z�C�༕�O���wR��`���X"�e5)f�e�_ߚ�_��M�	)+;Gt�Ѹ�6g���X��pUƫ7������eh�/�dO@Q4�$�U�@`,�0�g�{�Ė�(u��߿V��b�DZq<Ԉ*p��Ar���8E�����Ld���g|��տ�o:L�SR�R�?9mh����y��ѳ4�ŵ
�X��5�����������É���(���I9���c�gY��}�*��*B:�8��\Ƨ���H�F���!i�̺�Rb���P�|`�a9�
��DK�2�簢��%K4%*��A	��L&��hå􋗵T���6��qC�� � ,�L�
��J������+�}|RL�1���R�������� �k&���Ȉ���mP�ᛢ�F�*�h� 	�~G���5<�o�zƓyh*2���+n6%�(�v��Os"�:����{ɼ=���k����&����wn�@�O�E@�����3F�vF~$Qz��Y�C��u���4a0�_>q$E�E��##�^bʿ[�fp��j���uo9�a�����~*yy��<69�V���!�m�\��ː�N�r��)�cp�
�2硺���a�H􋱅�0�b	��3Ǉ�,�c�ojQ�_a���UP`Y�8������$f?}ͣ�ܿo��[�%����%�>3c^k쟻�
$�0a5q���e��.i�N�f�Ezp�B�|��	�]r�O�=:�$?57S2E/C�rq�B{>G�B�����e wIEE@]�a4�rU����kK�m|��DғQ���-��U�B���>�h��K�։�E��P��''f�IO��FB8%дϘ����Al�M8%��v��X�3��׃�������-���*�gs��/��%��5LL���p��p��T$���ߗQYdi2��:4tb�2눣�H=$��MW"0�����i5�X�,��ȶ�:��M�_J
���R櫙6�5#o��K뱄w:���G�������)��኏��yn}�k-ųW��3���W{�Ï6_K� |�����Y4&ni:<�,�"ě�5���j�@9U�g�O�S��S� �ύ��E�����Jd]�G��ѝ���>��k �fg�(�Wf����;�YJ��U���1S�Ǝ�b}��)�����)���]��X�P�;��T��B<���Tʏ��������6q� ��q_�3�'w����"���������6��"o��V�3���O������s���ع��𞖍�9M�<a�������&�"	�-���|��������H3�G2.����-��<�И񆔪�)�����-�m���x���y�mN$�gς:%�e��p�/Ҝ�Rcޫ�b��u:&������¸�ۧ
پ#�b�l��--�	<D6x��.E^(((�Pp�pc}��J���o����L�N~_����e�<�?0���;#�Z7OO�p#F��8'�$>�������M��A-~���uH����{�Pc����.&PE��9�����`ck+�:,���hd�YpQ�A��5p����&#M�������V!e_���YV����r�C		:�p��d���K i�093OS[�y�����B�̵=�Ĝ+�����*~6Zŋ����W�/e��y���)��t¥�qN�j!H�"|��r�DW�E�Eed�t)��4��I�8S$RY�M�-��&��B#�Y���:n�I�����;YP{1��zD+?���%F�9�pڱ�i"�<���@RjT gW�~��c:�{V�%��?�2v�U�+wŘmf��o������n�{,K�WW�<"C��ea�gf]��07/��8��j� p�&p��vYv�B�z�"��ee����f)U��^�8+�}�`}}����`}��S���n�"&Z%�#������rװ��J��݈{M�]�����}9�ސ'��E�7[׏P/Wʞ����9h�d����2uOh���,שHk''Wfe��rM�GGmm/lz��_�=�{�-i�TR�i"At;3e�EEnU����_5�KQ���w�;��_J�zQפ��MO
C,�k�Ȃ<���m��_&+r7<�Yc���^~':8/�M� A�o߹���� ��UfrR���d�$��q�l`��HZv��U�Z�8FO�hp$��u�c0�պ6ض�翋���"�F�̲R|���Fl������!�pr�c�:���5�Wȉ�����*�yuD��_��1GV�tum���j^��X����O�gCv���kR�lF�^<{��(�s� ���������zv��6)�� ;��6p��xa����l�O^JJJ�V��D�a���;���`�y.�������i�Mtܫ��Nf�������)>�vj�܊G=�� )0Αw��UU��&&�ߌTES)T��+!�C�����*-��jT��#�<L�*���)�Hez��� �<å���p�������N�R�g�E6�W�<HrrǟXXk �X*+�f���Rm���R���u/�2��tI��+�=�� �6����|a�&�71�+�!��KM?�����=��xz�u6���'1����tƏ׋�/Ʌn�Fp�.F�������C�D���%%ꁕ�e���ihh^��o�Պ{(|������ERXz&y�W_�"�����������%)�x9��Kr�QPϨ�i�3�扅�Ɋ�����5�ɯ�(��~��$INGNp^H��#&!���}��i6����DF..���g�(��S<'~wZ�����<���7O����4���+,�������T���3�&t@kt��.����1��M�M�N{����7�$δ�J�N�x��85?�.А��SKs�_����"��of��QSS��HX3k!��+$h���4�_o�ޏk<����<�3���<�	�R���!F^^�ف�4*h���m
��:�.�DHJ��%$������?Ń�D �c�^YAe�̵��&�4���r���5�E!Z�m��)�e����n���aLk����Y��[�3��ӧK(=6K�������kP�/����L~R���V�&���-�sr�*�0�k��t��N���(D]o��P&򛚺
z��I	^��r>��I�`3~�C�c0Nը���*��f�+}/�\�
��Y쑻���HAZ�3����j�BӃ3��(X�+<�gi!�z��Ċl�Q���u�ѥa����Su�JO��+J�#��m�r�8��j���� ґ]�Z��R�����������'�x#�]^�+��69>0 �IOjlmݲ%a���(�96&�cn�;M1�,{f++�%'���B���:_K�p^SV�3H/|�u|���xŞ�N��V�y��M���[L�L��Q�y4�EE���s���cb��y�6:�;�����}|��?p0s����X�&�J����=�lj�N�۷�9[�~�
而,���L�0��[�Bݼ>fO�&�<��J�V.���Y>�n��	/�=�r�)s���:�Oc#��oss<з��6Ų�N���fv����kA|��ڨ�ff����­������C��xD���M��jt���8_���P��nz )���?��w�ɓ:'ffhw�OQ"��>������,H��3���'�,P���,�g�cۦ>���=T�rt0�{���,@���iʐPă�\�JII���M���"���E}$�dʧT7��"���b�s��|E��g��D�C�k$n�9���a��S˘&�����)�7٤�Y����{{�)\��o%Ì���R���=ill�����\��6	�C��	�q�rDF2�-(%m��[Ȁb�=ST\�Z~�n��Y�%!a(�Zy�B���R����;	u6z��n��@��X9$�n2�����^�z�(R��3�*mx��(��\��?ҙ�oXm#8c�Z�l*�	Z9���f/�H�B߇���q��ȭ �����L��
B�R �J�L��ՠ2��ui����ћ��<���������z�:��I���٨#-�t�0��{-vB��/�B_�v\��'o�_���O������F�*�P��%�v�N_	D�� *�l���*�O���/����9�5�4Zt��;�{�VR�,��lZ\�`x��x�FQ���s��*�r�O��t\�5)!Ư�(������<�:�p*����Uف��?t(z�[P��.�O�-���R��`�vBa$n���6͸��v���+/͌������[g�Lx	>��y��FA�����k�����rvKNⶕ�������zI�&AV#w�S�����CK�s��H��",/Y�@#�a���ڃ�s�� ,�Z@X0��>Y ���B�)1Y��"V�;���w K%3�Og����w�_��q7�; =H����1�/8�wY��`z�E��|�J�t��8�=����n�11UG��݇ ��=�����~�0߆c��#�m��uL�z\�q�(��"�P� �olj��0��+)+�J%32��T��(����-V�`j�[卋=��4�.5�Ԥ�tC�Vh�TU݀�{#�|�uйL��e��Op���E��B�c�d��^Bn=�*�`@�����g|��'*6m깭�����> 9Mg"�_@%ي�d`��`�F���3�?������IW��Hj=z҂�D�p!K���
D�\."g��j`@��ޗov�f��~�>��T���%��JRg�.�U*��͕K(�?f�9�{b��@z06����M�.��K��O�Ѕ^E·P��A�AZ��4���8w.fe�_e�A�J� 2��Йc�7N]�y�� ���U�<i���nbHP���%��|��C�؊��y�!	�_�F�pM�i�aŭ�w�^(��#�?ۆf�s	$�6�'��A�,��/��-�Q�p�9-(8� #U�e�������oz��=�f��7a�_K_������?QXߐqcm�^M���Io�Z�p/��$��]R�� xV���w����>c�6�AM�5�bi���FE��40��Zx�	).�|0����ܜ:�o�^�_j�=����c������׌�����9
�x�~�
K��{11�̔����g"M���(���Ln�9�Mc�~Kg�<&��Wc����������{)��B����OMx�e-LpuC�8 H�:e}9�|��Y��}� ��!����W��}��P���s�"��+�U�E���
.�K��)����_�6,Z8[����_���U �&��[�5���GVS�o5���/��n���x)���;'g˴C��������o�QxX�e���������,�����b� g^^��	`�I%�~������,�_��sml�d�eO�cض�\n����w!]ݩ.D�~��I�q�:�L4�^��n���H&]^'Z5I�1?R ;���4 ױo��֊�.'Ϭ���G�]���b�{����ͤ[C���n�B>Ͱ��r'�z���G�H0��&+�΢�x���٨_�eC޾=�I�.�磕��]k��|����ܵ���f�-`+߱�X�_++����Ty�M����6ge��lnz0 ���b��Â��=FE!'"��ڤ���<����TŃiPc�,��롕�pʑC�����!3
Z	6��^��Ky���&d�O[G\�s:^{N��a�lY��@�^�"+?Y�*�F�]SF��o��Uy�(�Q�H���o������^M�n�S2,�����w�l�9�n�k���ײ��w�";��ؤ�B���]��5	|Ԋ�G�}���e��.CV!�%�x��#�<���%���b�nP*�d$-;��c�����bg� ��׷�������C������:cp�z�<�����Fl�C������!,*�C�҂�	B;��`��)+�I�_�g<�z�_W58��Ç�k���w��jZ�n氞���<j�����OP�e����E�����h��p��m�$�H��-1~�������n����Ai�r����E��.��ۯ���sd�m���c���������H@^�`�MP���W3�K�:Ս\�S$�S��SPxc��h�
0P�Q�c��;�!òq�ab ���	��h�ar�������>��b�:#)a��p�c����e�,�ۮ�����''��E�(��;&���#�z��:�d%X�
����8�٧�'9ȉ���/Ȟb��]Uf��qQ�SyCHpT���
�Wk�G��u��ō+�!��u�Qnb�/p���#�A{��4���)�������<99��О�(D�-�s,�FR���+�x�����>�A<w�Aĝ]�,+��q&�2(�X�6��-��.^��x���:^43��%ӯ�]��:3C�l\��g��E�[��N�Җ�9;��)�����ÇLADp�mN�e�����%(�y۸cH0,V�h���M[n�բv�a{+��g{���שiii�"r�Oq��_�@���|hll3?�؈���f�����ψ�l9�F��������������/�yT;�t��EE,�����O�-�B^J�Q.> ������gx�3�J�����}����
��.Xw4fiB�bJih=��z�2���h�O���nBa��o4��?�a��Ɏ9�r/�{���/���z�!߀KKE��v��/���ǧ�	�RHT�iƅɃ��wf�Z{��ub]���xO��QZ�Hx���z��m���5���
��vřI��˽σə.R}J�oB�"�O�59����f���x�Y��*�1]�r�HBB��K���*�b}��i��i]e�jӨw�Q�K�^��O#s��w���U�:��yǆFqr���(�G��%��lB����hV'�$j�0!A+<�qUkѬ����嫸���Ĕ�����f����JW��򔒞2,u|||�>}�[���,]N߄�>����d(ѓq�7b��}}=<��95����~���ͽ�Fu�d��ޭ�t{����G_�-<n���̲�?��8�חUe�m:���XUUPX�I�{be$,<���7�3�x7�`�G�2�_�\���B0>
�C���$
%
W|Դ�q|t���VA^���#'�ؿi0��CXD�ҎM����^[�M}�e9mtd���Zr׫�~��[��ܹCKC��{t��UX��ܯ_�Ϟ]4-��&Z|ŀ�$��������@.��4���]�|y�,�ԤG=wk��*>��Ϡc�$--o
���*�^?y��cs����nAX觭�[�����Og��w�ccMk�<g�+��8���XZO�Pf7�F�P�K��4_�i�/ڞF����0��lȷק	��989y�\�$��Z�֭2ڋ�M󲲮Z��pRX�qg���n��[2�������ٳ�j��h5���x�吿677���,�udb����j>�� �7;�Q��N��p��o o�jaaa���IS��6>A�\��H�������HZF⦲_B�:*��N`������)mos�H_��:;����/��1��@����� 2{��˃����.v���I����D����d̠1�Ztt��<�4�	���������)#P�%��
:�J� �BCm.�='�Vx8:�7������ѨD��!n�;KLOkkM���򴆆���\o�e����u_]Aޥ	�0_X��ţ�>S��3M�0��.������P�������z۾V��(��J�O(�D����{�g�x4s�s��b-��g�߳�$zAp��qB����=j{�>�����L��D-��jt��pr��-~�x�r!�38������������Jm�_�n�*�ȘL\�7M�ѯ�(������m�<�e%��0A�fMNR��E�KaW�n���>\���_�H��L�:�B�s(��Pn�Z�I���tQ+��M��柩_�Z�M��t�k����on~aUWi��:kni�*-D"G ʐc�;�ijJ��ۣm�tG����prv9�D8�������?��>EH��V�F��2K���*�f�^ΨsO�wNI�d��J�u��Z|<�;����)hp3�[P���ټ�[衡�	b�=���h�O��iR�^�=�
��	v+mMty�w����ei���g�f����bi����z��oB3`>n�����`�%6�ʍ���@0��d���P>�C�ml���6Qh����v��-�҂�������[)ii7�;f�Gl������_5Sq��m�]�{���%��ޛu�==ʘ�iY�D-	&n�Z넆���?��-��p_������P�[y:
F6L{�*O���sh��`ajǽ�L�v�P>%%E�� �����^����d�~��O+g�����8�郛/�'J0e��݅�?��ƣ;�~7�1�+���}Q�=�C��jt|��k�{�������3с_�<�����͵���'%��[�m3��y�oݔd�ʏh����G*(�ڑ-+s�c��?��t=,��g�:��A�B��ɚ ������^��:�P[��z���Z�v�+;55W�����c&n�LQ�� J��Л���3�$2����Պ�1X,�Ma���W5M˴@���@�6��~*��ө�h�x���D��bʪ�KR�Y���z'��	H��s�M6^����֖��\!{Am|L����������O�蒐�X����_��o���D�gQj�j�� N��M�[�S�c�8�`|��ring��?��ݿ���L5� �53{���M�a���k[_5r|9BQ��E�X9tq񣃃����.Rny��c\�]7�N�Q�gR[�yW�lY�������#P���ng��\���v>�)����+U�f��
Ϟ%d�8�f����޾=0?�����'Կj�LUG�u�������������-�9�c��}$���O��.�v{�!�K��/loG�G�c���
��+�-]\[Z��sPٔ74�ttt0�L���+�ݏ���?^u�hnP�T�,�����B:!�j��R��������
妧�� �]3rMR��|b��[S�a^K�kk�o��&-�������4mu/��SM��u�
e�{�Y�\�A�;�GE"ˬ��VE���Tء�.����< �,a�蛿���7sww>7�����:��|�}t􎶦�0o�ewwwEC��z'B���\�^.I!i��[d�N|��ޞܮWj�7�,Ĩ�9@�����^�6��ֽ��<t[����p�*u���[Y8����_��>7q�"�ry\��1��=F�<���O�b0��yk�g�t����*J��ܤ������>Yl�v�7Gu�����r�1�CV��1˞$���_�W&�3��w�����.]Rzwʧ�����*��Ν�b�s|�Ƿ��L�=9]otO�����?%J;�x4<�ZpY�Ҝ����uGh�ڏ�o��ߛ�
��e���ki�g����8��N�=޹�QZ^���:��~�]/����u��FHHI͝�����@�۾4+��誷����j
G|9�>��t��x�#
�4��d#�9�V���ް;���:�34�xL�6�o``	��U���|�<����f~U�#�Z�̯!chǅ��������݇U��N���e���l�pq�tT 	��j��WA�m.��tu��n~#�l����]����30�|1�N�9��a/`�@�A�g���ٹu���k��;;9��֮��>B�{�vk�t��M���P�S�9�T����eQ�:>O�{ob�UD/�蘒��6�j4+��L����/-+�=3�;h}O8ݛ&0ci�&[�~~nN�w-�	ZYT� ��v]����*D�<K������#�<�JC�mv��ӲoO���z9y���=��oz��-�����mm-}}#�n����R��޿%�Փ�Eu�w\0Ԏ՝b��v�h��f����W�����e,��~�>7��d5�L��8�#p ��D��N��~c��v�����>>`
E`Y��� &��E�UU�vv�C2��H:J��6�+�*�Ch���:�����EE6�</e���h�e��:���������w�3��i_��˙zv�p4�o���v����o~��d��!ꕝ}M+N��륿<�������<@�aw7ak�e�'���X�i.��J�d�'��}��T�Yj�����.k�YC[��z��_<�� ���xl�4��II���ISB�,>z$}���Tέ�'��^Pp
�H�>y9���ޜe�c���]u�dT-*�urO�LOgsrq�(?�/���f����Y"ş߿���p���tvv������x�V��/^������8[.;�![�>Ꚃ���v��"�[.�����\7���̀��uO��2""��-ncG6b���C���,�b��� ½�ի�����F.��B[u�<c�lml�XG����`J�_��I�2�!����݆��[$[��-���w����f�W���[����/���{���D@P���4��~Q]�Ս�'tttFۜ(�|		����uH�FD��9�O�������*��>3��c��oΤ�{�)�q���Tv�KK� m�F��D��2F6�^�g#g��<�=�Q`�*}N0����ښ����z�O�}S��/�VP�od�آd��ַu�{��z�mQ�6�B���Z~2��QM�; X����e?8��zz{u676����M��:��!V�����6 ���?���`�L���W2+�Kl�\l\t[�����`c-��~~Ǩ$�u�A#C�̎W�Y�����nL�j){��&x
���;����E.�mP�k1z�b���4�lԡir�U1cg^�	�l�6s�����������z�uʔ���ط��ֽv�f�I�n߮A�ʋ��z733�?��=�s�{���@
��� ��)����b�HW5g/r|m��t���O����:Eʔ�8���*|W�6HDŞ��������?}q9���&*���C�c}�%�ݷ�&bZ6���s����#����s�0ߜo:wLT����Y�^���2ۘ�2+Pc3�[�)c�}S���l|R�[y>������N�
����m��v����:5࠻���l�N
Ed!k)9�Bv>>E�����ʷ������z�t1������(�!Dun��fB_�w������b�R��ۗ扻���W_�<��N(�յ�?4��=G�V)�M����7'"b��L�3���|*�y{�u�,-E��n-�p��X�������:e����ߝ�FGF�4ٽ�|��^TП�Eu}؊�M���Q���iW�ieH3Z�����Cչ�i�c<�Nnb4??�Az[ |��M~@	� �[������ŧC[3��-χ��G��1::���j�V����nj*k���5�0��11�4GD�]��G��Ć"�Y�%h;��{]}31+����?��������4�i�Bh닻>��nm݋9���ɛ�ϩ�[��f��#�ml��lwhk�\�Q��d��h��Лԡ޻��"oІ�J�{���,������9y{�_����,�l�:��8Hp?��^oqii�1��b`45��@?�S��}�^���	/j��6��p2�����M�+���BU��Y���«S0�;���Hl�1O�Y͵&�Cu�$���
��ؤk����Z�qi;������|h�
7�V
�Ā%@|8ڪ�P`Ѱ�}�ַ�>[�:g��}����ʬuz�6Om����3���K�D���n���N�KIK=}6?d?}svvU���l5�`�I3�>�
�ʚ���/���:,�>�1�t�����B�:�pkfx�=x��iu#�nm���:^��pB�u�0�hbR������sxk��ϝP�B�����υt=S�8�߆�W�WG���Ū������Δ̞|%��J"�T����x���v����.ӭ�QA���[�@ ��c�w_D􍜤��{`��xs?"��k8���\���d�a|�5���s���X��  ��,O�!~��G��M�d=Ī���`S����}�R�m�,Fn�g��x9���SO�)��f>�t��4�ql]�kae����s&�J��0����
Ň7�{�5�7RM���.JK���v?7z%A[Q"b�=�$SU�o��K�?�r�l{���.��H�/���N*���W�F���x?�8#*���8F�&.nl`E�y���뷧��{���Ò��������G�0�-,`�MdJ�i��Qzw�A��aPH�����K�>�/_jI��ha�ﲮf�>���33#�}fB��*��W�÷�o������q�	���;�f�>.��M).���Ǝ�x��0 ����j��a�&�|Mv���>��*��OPK=����c�ӂ~%TV
����G̗��=*�L��Tp�CX���9�ow��O�[��ȚJ�	��z9D]~>pr�����fJL�@&_���1��P�{^�q�(��w_O�J���_�<����&�sa|yj�0�W�Q��a�ٚ����J�?�@�WkiG^r��VXK�ﻶp�h���1��UP��]�S�o<�0l��<�:t,+`S��׍r��Y��`Oԏ��d�6�$�!��sX��iqp5o��Ȑ�]j�v�dis�$`�K�4�t����eͼ�M�qw��侙uo���-bճg��^������p�I"�90H��Ν�tAa ��ը�*�|�IO2�%�ѱ���}0�K�Shl��@?/�����֝e�,F��������{ݍ>:*G��� ����[^4=�P��U���d%z��5��@/TBˠ �����%)L�d��M�lt� =���w�2?�̈&$1VƩRX+,�a��<6E߶{�h�
GG�ӚnN�|�`��`�H�F�(F�����J���o/;9�����a]��7W�#�������JC��W�C��D�����_��%��=f����D�M��>���:F\�r����]� 7�\�v���r���sЫ�;��*�#����y��U�UU���"???�63�lYK˛�c(K�����?|��ԣi扄���=VTU��ؠqw�o��~:�-c��b����6�������!��k+�4�h3�|7�M�C����,����5��l��C���I���J��ɼ�|k�}0�6N%L���i��\����L���P����7���ia���Ðe t�����-�O�(/P�8p�6,�t����[�D)Q}���*��ޤ�3n�>�]]7.E��yg(��ڒ6��uV$�����U:��z��lPx��כ �Q��Հ/���c���O-|�v�4~�݉�a����N�W_��!�ܹ����?v��)�M͂7�Y��1��R�:%�~�S�}˴î-��PK�qW}��B�p��nS:�� �=8���%`yP�{�d�� �vb���X���{Ga���$��d��ՈG2KY����h�Q�ȯ����uQ��؎�0�l�c;L�[>R����=ZM���|�L{�=��յ�����x>���&I���f"�����vgwR��I���曒YV+XVA�Ap�F��SB���G�q�5��z~I���뜺L��À��1G�%000__�3MDOo��-��w{zEEs'>����p,BZ_���3OL{�T3��5%�J��!�����:��E>{y_��`H\G[5�>"Q��h�{��!/�l��w�n��}\�嚱���k8e�Z��Ύ���忥�+�U"���

0��q���zv��(:J#��c?o%"}��[����>�`Et����u=+^�����1_jO��D_O��LF
7~A��}�'��fDDFV��+O;�t͡&�i T�r��LӉ��V�gCv�pՉ3��+�펙u_�^�<��W٭��T�T�J�7qŨ��)_^P�����L����<)׷��M��R�\�������)' ,`�^��&�T�N���B��8�1nK���,ů�Cs!Qp�a�K���Q�6gL 
���VA8��g7}�����Ľ�:�5�bdp��-;*n�ɶ��ib�}o��P�q��|���`����W�*��>2��8�~�E�a�q�+�+�ݣ�_�����7m�w�Y�O����A���I�iy*BuFpxlL��Q{��MV��d䅔�T��Tm8����R&3J-��N���VaD�@WwwEU��2���:{�{��8q˄�~�}� ���G|���^lb%C׬���a=�y��I�++���B$�H������<�g0��R����h���uT�|����FZ��b۷����E�0?V����r�no[$���SH�ˊ�����s6tZ������x�K��>>��='}��

nn7�b�Ġ�����������[
뗉^U���6O�X�cŮP�����Z�_�
�ۜl'��v����7�~�!��:K�I�"�!KsF�7t��..9��=q�G>Պ߿A;]�&u�E�Ҳ�����g�Oy�^���0����zA�t�t�}�����L�?
5��AJZZ�f�%2�� ��j��e�7ݳ��)وL�߆����΄W�=�����8+++�X���`����G+77	d'������)C�?++�����M�,E��~̓�V�.���o`���U��u�^�Q7p���������Q�k浇˾�/e����Xp�	��P *M�M���>��^��[lS�SBO"��	���L��3�O�:aa������:---�	T��~��g�&�9� �'�q�-*Z�y( ��O�o�R-'!%������f��8�c�4����c:>y�A�G�����e�
a"T�!ST��G������A]==s�]S�~p����{{{��" ���2@��;�\`����:vj��ҡ�pq=�ڜ����Bo+?{�c�P���q��9$L.W�Ȝ�g�Y���Wou�������Ւ--��(Ym�e!��,c��F����졲�J�&T���(d�R�&&��3s?��������ݯs���z/׹�G^O���sD���9��E�.�*�O�3\�V��j��Մ���历_�UQ���K���+��V��������ˎ,{���_=��E�/�QTT_YY��Rl�Pﳼ�jv)x?����D1�~�/�W*Y\<���7%����22�~�2����4����'Ѿ
���0�&��9�2�߅���-3M���]z�)�]V{3'�{{꫰��-Y�9��ⶀJ��K�.��R鶰��r�2 T�^��	}���k���� 9>����a�O]ll����A���ꔕy%�����_��[�{���Xp� ,��t�S�2y�-���,��]ua���}�m�����r�b<��B�{��Tx�W�_�q))))��w�}Ꝭ�m`�+W��}9^SS����C�g�����|~{;*+����|����?:%�+vra����T!#&JO��������
H��
�ujW�*]�P��+�Y2�p�.}~^9����73���0�qQ�"��ߔ��|�/E,���'���c���=����A7;�+m�I����"��::��{S��K���k:�(^��+���U��4|��S�@���:�;^7�����p��>qږim�{Ğs�Xj�aƥ����ɫ��I����Kbmdd�Y��`��������hЮ<�oh�������5O������?bt]�,LP����q��k�+�]�2	��rͣ= u�!���ӝ��,i�M������
�v��y�i��޸Z��ձ5�HH��-.$�z�3o	*�E X���.�������Ӄ�怷�#T(�**Y��K��꒢�֙��vZ��� QN�������}��?�޶�6���ގ�Ћw���KAA��ӳ�/��MLL��[���q��2��銊�#C�N���nh��\"��{�fq��1i��;-������͵SE�Q������O�������_^W�"'��[ZjUj�p�MѨ����f��yiiihK�b=$Q��H��
�DM3s�?�72!c���'��2ԗ��@|���OmҸ�066l�5%���f�Bw���e+���5qў|g&= µ5�?XKѡP(��5�o�!�����ymx�p��l$�Ç�FG�8��GG/�$ܸ���V�d�z��ŧ ��b��*�"�Κ;��;Y$r�n�s��#�����z��ŋw��U׉%�u�%z�&|���;32�]3��6�[d��CX#��D$H�۷o���.�+�,����;Z��(P�wv��Z�5���ɯ_� jÂ_�|��5�p�۷m�&Qs�*��<73CJ�=��4�ɨ�S}�߭}!))�� �o�Q�}��1�Sh�o�^�ݽ������Ҿ``o'?�3�a	��?��e��l-v0]���|�Ȧ��@x
N(�!��v�`X������
>![�}=:%���nm}xK��L&������L�=�������	���Nb8����Ƈ���3�Vig��qx������,0�

�CC�0Ň���A����E?C�.�з��|�&s&�����D�=B1��4{��s�LDf9X?:�<�/��h��t��@j�0�,�iei_��終ώ�<���Ó'������M�|��u��09�ap��	Ԣ<��87�����G�\R�UQ]]ޔ�'��hk;�Yk=V��NGG��ԛ�R8�����@�������� �[s�G!�Ү�@F�FrF���!��x��7T���ҩ_� �=L��!z����V��I�^Z2xQPV�>�U8.s�n�ؾ��0�ea��O��+�k��]�|ܺ�r��M�ߥ��Ӱ���w��"�t۸O���M��C�2��
�k���(ͨ:������V��`p�"�_Ł�{�Aw]��vq��}.q��e/�`��,oHw�X�M �f���1v}HU�zWV2�lٲc���	��))�9D�bEE�#5�K}��Ve��Ь_@J���ˬ}n�"-b��vf)R��)5F�W�Ė𻜪�T�t����__Z^���Br�Qi��c�kA�����h��

K>k�R���atj!#�4q��!9ע��J�By,�|�=��x�&
����Ԕ�W��J���J���[��S^GmB���h�]����Ꙓ��{���©���:��~������������쑻��`R�{Ǩ���@��S�ڟ���li���R::n��t`�c�� �Tq����]���&k�Vʘô��ZYY1nsb�h�/�#��`>'k��+"ӿ���o�){[Ў�!<TH�s�����)W\W���n,�ݘW�=�V=H@��S2,��	� �<�L1���AKED�uu�u�����q2)D[V��O/L��t6����EG�J�j����{D�^��KJv�)w�L�0�4j3O޵�*��Y(S�{��;:���ז������6�6�B`��jk�z�vlD}*���#�-
Y�f�=C?@����uk� �\+�L��C4;�U�6`_���65|���!�w
��Q1w8��{(D�b�L�T���[�0LQv�� |�!e��5c6��t�4�5���yy=Q��Hyd�<�߭T^����7���5s��^p��|��D��kW<�:���p��UL��O��~����穽;7�C�D"m�\��J�E����d�ě��~z��L�4�ş�����ǌ�|�߈�SZ��yә ��Tb����@S��]�9�W�Rk��WU/0��4鉠pɕ�G�w�|�j��/��:(0���̚�qg�g��g�m7�a��X�%�5ƵĞ�ޔ�?i��&󨝡Lˏ�y�v�)�@r������5Sy*������<<�?���}�f�/��Z�����ξ.��;�@�?T���n������y
f�/�eW������g�m��K�C�>.++C���С����������ʸ��6%���d�t����P���jo=$�h���=F��X%_��1Q=~&����a�������k�d�`.6U�^d���ݎ�svt<������TESS��ݷX���+`bll���+e<K��ikw@J��\��G�@vddCj�+�Ϡ�g�Ev1�t^�"��j�ݨ.�Շׯ�AG��=MJ�(GT'�����>���s	�		����$n���`�+�3X^^���7\H8^�����,wQ��@�#:W����ݭ�<�;��\^�����ޓYz���J[�K].��B�Đ��/J5�L6i�.7O_����K8���Ŀ>;/"�J-a�A�}�Bz�ϴ����Ctt��W�u����=�A bl��ӂ!�]��@>�U���!A����)������1�}6{LZ:�'�i�a˵Hc/���B@x���g��<�e�W�d�V�}�n����_�E��ߌ�p���FAnL��!?�=1���$:.�#��^�{К[,�}bb�Drr2D<�$�fvv���t��HN��ڝ�||�R2ݻg�� |;6�t��7�fm�XF�쬀�nW������� X�o��c2j^qB=�sq��<Wa����������r��q[*jj�XXtoڙ�^�	G��%�%v�"�������>H�������+���5��MMi�~ yq8��dgg����±b�.jycc!�H|�.�D��{�d]˗P�@
**�4y��s��^f�F����J�v�i�s�U��Ó7Ng.8�SVV�+F`ejzA��%e�0��b�d���-,-�&&�d��/���H���� |,l
{�C����	��wM��?���tO���6E�]��	c����O����V����O$��~k(-z�[÷�e�	�y;��o7uD�[�=b��fV�<�'P�B�Y�Q8��������������ń��/ttt|����.&{��,.���xT�~(�}G��}!�*G�Z;���)*�d7>a��oĕ��E���̻*?��P%G2[� �-ZP1��}t��E�I�A�D�-�Ʌ���#������d�=�aO\�aXX��̔O�^��ȫ���^	����;�NM�*�`�r�n�gd譴&$����)"MAV9Y~�� ��_��"-�����\�<�ڂ�a)hz��)�LFG���SDFN��sDD�ĸ�qEg�V�թ�隁 >}����w��<o<�������z�������6sPt\���$��X�剠=��L��_�jt�>Ä�K�;s�L���d�,lXEʃ���E6��uu����M�#�[�����L }J#^���8�rkhA�ð�N� �z?[�q���

f����5��o�?�:�se�kj�b)O)�I'����$�jӹ����J�[���D-��>)��7�#����t��&?F�ۭ��r�9����W;���q�������,r� �9����skFx��I���/��5,M�
���LO����ֿ�Y������� 9Y٧���)���T [*՛_@@4�!�p��T:rĜڥ�诗�)!?r���VVBo��F uAt v~f���E|�^MZ��3>o2��8	wx�P�腀�]؇^t��$���l��5��8�dť��@||��ܻ�x��w�2����h�����ݳ��J���[�5�z''ol��0K��|t���jˆ���ٌ�ޚ���#;���1�SS��q��ZG�3�**v����nn����̨D:�Y?�ևd����0��\-D��]�#�f��\K����XU%rcC��$.G_Qe��	�_����m}��5^n��E�xo6���G�Ch���z���Գ�M���::;�_<M����7JԬAz�ZAa[jZZ)�D�ڜ;������heȆ�mш�+��C�.��m���fF� �k��'������ͨ��sX�7�5�y���߾��vC���O,�0ͼ��:L��\�q?7�!�H��������6��:��5��J$t��W�ъA���F�r���o�v9�����J$&0n_IU��ř�!�'���LH[�D�XI�|ӦR�Tb�{yUU����jH�e4���*�tJ��qb|�
��WS.n�=59�T���9C+$��� |��a?�`
0 �D$�[u�-�2���P��Ӎ�Oʹ2ܷ�	�korj٥	8�~�bOb�^�����N��j��G��J>�%�����ڇ�w�UgeYC��ޝx:]C{����nU�n,<Y4��'x��llc���,,�@�>!MHެ�����r� ���͑�ԓ����岪�� �@�����n���Z�;I�]td��1��ە��8��i�����埓�Ew���3WH�_?F��)z
�~��������G��
��/xB�u�n̿�w޿m!�W�����)馼/@/���ܕꔚ��A7�+\ve�Z��C$yAډ�cJq;l$��3%*=G73�;��"� �	�jɐ��)�����#��tB�����l��]s?kj�	d� �A�W�N��,`��D�@�E����Vk��p�"���I�7T�WL��?U[��t�����=����'�v=��u�|��>`�9�H+{�z��^G����Js�4Nt�څcF�>�z�x@�3@����h���!y��v�����o ^Ss���QAQq:t�y�y���
��:~nYi.|`&d�E��BC1���J7{{cF7u�8��b�yA$\��G����,�6���Y^F@���<r:���(s	�����5)��,҇������Nn�k����2���V`H!e`�w�И
}7a��1�f�Sp##6VV=�O� ����|��,++nh���c@fQr��T��׮�G��i+�?��{V����i�t]���Jim��ٹ������7�9!~�RߠB6�ÚC��sO>޸��Ѧ���������z�({㶤{k�Xo:�6��7$��ܢ2�A����{O��$��-a9X�BJ��h;R:GwA�0������P3I3�x��rN�;��gf�7]g:A��`r���]J���_2\co�599�d$V�����Oo=_6��p�v�����/I�\޾��ƙo�jPaֳ��M��>pxG���d�\��1;��Х��ߜ�XN��\�066�;l\;XRY�bĹ֪�S���=wA*����W��oE�*3�}����r��4�$50#�o�Ĥ�z�/9 �c^�`Z�	ߙ�zQW�<�����RJII�0E�&���H����V�-z�O��L݀4ٱ6tt�j\����۠rf`�Zh~avP����K�pkg1�D<���~��ZQT���%���gYJ#�ޱ%Ŏ�o�j+rC�.n}��ME6lx���{�S�AV	�]-'�uSN��Oт�F��ԏ�)%d{�6t�a�	v���L%����'��)��C���r㢽�������s�4���KP��2�y��qE8���DF�Ȭ��^���w��?�V@r<P��`�*~c(��N���]�P�Ha���Z��ZG�i���u��l_[	�eb�0�D��c|ㅖ�E����Ś�L�
,�ȹ�Y Ƛ�"����p���q�s�"�g��!��cW���P��d-kC ҿgOk�D���������~~��IZ�Yu,`�v[�,1F������2�6�u�̟Ǖܻ��:��B\�Br��I�G��ϮW:�2�󖽽D8,,�Z�F!���׸n��+�i쁥�-�(Q��� }ĭ�4] �[���z�V�%w�Rː�Z��l\*����kᓱ��g����96�|�%����ŏ6X<�E���l�/�]-+sY��Z>oh�*O[φ���kR������ʪ����=�X32.���+�M��*ͫ�2+ޓΆI�ɤ����L�� Za��W�����f�10�P^�P���s�E�U����ʔ�e~!���a�Ɯ�!���k��9g���̔��5Ct�(��Ҹ ���[Nf��=_��Í�6]Q�"���#UC�huMv%e��(�Q��-���Y�w>*�B����Srs�C͢N^�:�?VfY�g6cX�����=7w����Ϳ��F�
�K���ۂE��rso�������77�k��L��1����L)��]�h��7�C��o�ml�7����O��p���9�fiQb����v�.ګ�`"�h7�}�&�&z����75S��<:�a����>�7[�����|�5Kˍ���Z�m�S>�.2� 5t7ĻU�������\f��K:v�chu\P@�}MC@>���׶��dz�����0�+����+gV	��0�W�mҸC��Nx��]�^�����.��^&�u�Ndۍ��b�8�@t/;*"� B@����i��g�b�=u�w2P�N�Wl�tK�\YQ[���DY'�S�rqp8c�v0 SR��v���&��gx���Rj;=6M��6�`��1#�0�q&j�F�rei4�Ce�C���(����Ak*�̦�Q�_�}��Z��C���6+���bî��%?�h���>+L�ܔO!i��Aw�s T�8��X)���_Dݚ��n��N���3S�!���:�hr�mr^���O2��͘6�,��~�X�y;Gkk5���3V�.Mt����z`�>f`�s���X7)}�^�	�4 =����P��)9T��gJ��U���֞�!�S��t	UCh�e�n*����E&���u���3ƝƋ����E}�a�j
ƶFi�߭�������V�f�Я;7`φ^I������wz�T�o���?�5_<�o��E/G&hΦE���G0�C��ֹ��e`^y�2K��":��q5�����\��:5�n�5�@��1/�wc�rr��_��q6���]+==R���{�ď[n��NMJJN����h�^=��<��2Ǳ������C{��q�}2�m�r-���ʦ���T٫�cHe�m�+w�k�0��#0���7n�)J���3�*���;8�F-"Ħs���r/o����hȭ��.����~N[w<���>a�6��)io��I2*%�C-�#4��w����l��j�@ ���-&{j{޳�[�qnra��bߘ|真��C�J�1�ƛOi!��7���F]\\D�q�W�)us�ҞI��;[��p-z��0�C}�D����IY@�����M疖�����8�2S���r��i��=��8�D }�T�פ U������;ZVV��\��se�:�A`����<�>�M�V$�-������"_*���}B�@Ƭ@�!�vG�$j:ySo�~j��q���ő��+�l��.��HOTe���+ �c�����aG���u�a%��u}����믕�S��B�DE7��I�'��.]
�pJ��A��r��$v��W�SqII�t~����/3@�[8�S |��0\�M��*|�n�J�cY���.�`�ii� �_^~�Xp�ā�5V]�ڰj����uto}�|y��[TjG��TZmm�>��U	,��ELh"aLV.�@29aD~�bX�`�b �]�6��e�:��P��y��ϕ0�@�ܜ��񮾚�ӻ�m�ҧ��{񌾝g76 �p�ڥ.s���;�ZfV�a����lR^^�����b��d�9C0��kj.��RK�K=��i�ZQ�����WKU�.��E��/$��LT��/��~"+�B��Z@/�8��[�JKKKM}K��㓟�^5���9�^�m���O����v���U��S폱G��ۻ��sF]S���4�4ݹ�.�Q(F2Zt��Op�%)�Xi��kf[й�v�E	�@�Rף�����ܫ�Y�C�=�u�N�1�
�K�4�AG.4-'�!�zN�88��?�dK�~Jȇ\\�Q�o��`���3>|�&n�����s"CxLsi�Do���`��E'ｉ�}�d;���|����	���J;�'�!*QG�l��������Հ���Fy�S;�uܧm� Ϙ�u�4��= R&��{�%�WF����&)ɫ������e韸��S�v��U���ң��. ��<��3p�x��5] �\�|�6��D�iiy�؅�mQ��wv��u�$��qT�K��A�q�%���?��y���08G�(SwZ믤����!@|���b1T�;?P3N��K��9��1��S܊C�xMmu�����
��q,J�5J��6��Ӛ��q��;q7�hGSN�r��&\��'���4��^&1ݵظ�v�y67#��r&�{�P�m����ڔ7u�u����l1Ցv�����C�.������1~�/�:$�*<�FY��d��k����g�v���>|���,V��<G���7�5& i�j��8�-�}��ݘ�Bc_����iŝ,������ݗT�}�0$����^<�Z�x �8Chp�0(Ez�9�,�h+�ZLzH,�fo���Z���;WVyP�����v`��#���R ��VK6]���w�0��u.�q���� 	oC`�{�f�$!������<���twOO"D��l'Q���c,��!��`[a�9�.���:�1ݘy�dB����&$���RrM7G\>�-��]�g���}��f�����x^�S�X�*���=lڷ�������d���ʚ�/$`BL� ��>��J��,1+>_av��l��זa�'S�?9 "�q�\�`�fk�A�z�Y��,/
�1��q��;�����UU/�	
���h<��4����6W�A�'|��]�D��`�7R�b��&h����x�L[n���g���j���]}�"�����*@7�����>���4��:�Jd7��n������
ћkl�젛z�Tk���i!۶�����K���;�x�U
��M�$����7.%��(J�C\�i�Fu�����c��%���܍nd�d��-���d�[�G�Ú�HOc�Ʉ1�R�>��jm�ҴB�	���Xp"�ԧ�Wt��r��Ҧ�A�����E=�E����9�d��������r|���$/���ri\0iH��{;��o������C4��<�Ǹ(gf�\����2��w��V�Q��
khr�6n� @J���k`���r'AX�@��I�9?�O�YZz)R|�w���Gx)Xt�'������(�$��E^�%"���[�U��9��[t+��F33c�:U�[潉}���ht϶5o�M�clB��4��_Z���}����kB�oO���O�-|�p�����y��l�{���}��@�6_�5rP�w"�5���99cl:֛���~Ϙo^�.o�T|�}J}R9-����g�R��G�:yԨ3M�XE^���s*��ey���l��s�M�=P�2(�/f�8H��ĭ�%��	0^� ����:���;��ew��˩����&��5�8h\��6#W������VC����La%�kgJn�+}hb��D���C332�<�'�~i�)��c�*e��(��=��X�^p�m��q�۱���5�� H+���>
W��V�O�������N&��}m�0|������4d��n`C�1����Ae.���q�2s:=�$ȭ�o�B�3�!r��3�w�A�,-R��Mpe��=�o�9���3ss���'�85ni�a
l�2��K�d��h�({[t����Ύ���E�@���^W�1�5������
�Y�by��rG;W��+$= �ܢ�XƩ��y�YX�x��죀zL&��U��͗_p����?�щ󀇰��q�\��<���������sv_h�t��>���,lP�q�D�S��8$���+���N��>x�;��A�AW{�]s��e����T���d��J�ߡ9��:�q�
�v|�����ƻ�A��S����6��Yw�:�ͦ���^  ڊ
|q�����׏291q�Ҏ����637'uJΊ�L}����F��ٿG�CW;� ��
�gE��P�V(���Wң���v@���	fffIN��كt!PV&���y{�-����2��`�
�3!��4z���!t%�r쟋IŶ2�5m�k˵�3�d~Y����yW�h������ҟ�h��F�sC3o�V��d4��5=�\�%Zsgٙ6���<O7|^��$�\�\F�(�d������d��Ø��O���~�T���}�f����Fx�};�����nP�D�@�M!v��s���/�kγ.��q�;��E�!��4��4�.�(���w9��'�Pҝ����#�s��<�:PL\�H,�A��L�o!��)ߺ�X��1����'g$�6�����M�g�%�wSb�'�~�V��o��
�u8�����lsj}�����G&�=��<A��-7G��`�ڗg(l^��.� .yqCa+}�y��q{�ν��ۿ-3$t�������A݌ǀ �V�;�K�ݭ~P�#��b~����w��_��,/��qQ�b�M2������<Ig^�Zp�`��lN2KZ�n�[�¤wf][��9��ZO��x�B=Qx�����q'��΀�hH���	P�Y����(�����Z-K������������;�*w%��TZ��m�u]�P��-�R��4�����i�����չc�k�ux~|]z�p�9p��۰����II���~y�����x#�5�e�v��qp#' �ε�*��`=<,\ȿu�2h�L'^���<um�^⋧� z���;b(�\��Xb(���?������S~�oqG�kٟ���:�+�˕�h�4��t�!�gȜ:�JYWCײ7�c��!t����D�8��uj���N�� �v���n�7�H�*;�U�0�� )ɮu�t�8	�_eG�bz%���S����㲣�N��|�B�b5e�ŏ�0���r�; jb����n��ә��Fe��
DY+6�ymϜ��	9���f�q`sD�I�u��AjzzO*�ȏG�`?~�����h���,J\P�Q4ں?�b;��&k	 kq��e�Ly,�Er���_	\��2)s�o2�����������_K�#�9�#�K���p���S���j$�<�y�:|�*���9KP��� �h���vU��׮ᓚkC�Q�?���J t������1�W.r]�^i�!B��oD$�ġC�\��Ls�T�n��U�e���� ��fN��E�V^�j�D��~�5V���&�����oZM4c����+A��>��)*Y����Ό&��0�X�V# A��|w�3�%@��Ж37��Iڂ�3o�֞�����y��Y�k�-�ί�P}rle�3O5|	����u���9끭,J� 8}}u���9G��(4.��!Ϥe�(7����?���J��Z��芠����:{����0�A`7�؉��B�Vu���H�Ufe��հ\��24s�;�xv�j�������o�)M�� \��]e.D�Y���,�Nf�iiğ?on����s:;��Ԕ�+�ڿ��x��������]��S�//�s���rϟ]�$��ӕ�����rU���	�4�ي�G��--��X��be����z�w�����o�fΧc�J��@�x /�$v:R�
�-l^��Ҡ{�b"v�!3�����o�����mm=��$6lW-YU*�Lh��ts�� �5`(�8㤩9��Z���@�}��� 
�Ʒ�A��!���wa�-�4�WwG�����]��g�7�Vڟgi�����!������!3C�!�ˡM]sb�^;�o17f�m���(�5Ue��V����V�n.�v@޼>�!}U�J�[Tw����G�Ywh�����4GF$yB�V����C9�aa� ���X�ΑN�^k���F��+�L+]��-���<���T��F�.�h ��|��>ey��1�ԑ#;���5U�3-K��cϵHߒރ��A���Y�'���++-�H�C���3M�C��ۏ̪�qO�����
a����m�7^݁Ef"SYE�y�B�O��i��ο/�X��5�?��c�wÚ�-58�Z�B��E�t��`Q�
�vʗ���N��fo�\{����ǆb�! $���D1��,�.r@a��A��d�|�zUI�[�Z����^����1���[�{�K�5�������]���A0=����f�W��J�3�I��ip�-�]�.���d�RZ�R��j���FQ��k���u��ČP��T%K����z��\�DS�h�-�ٛk1??w��Ѵۊ�>��AyT*���M����S�����<5N��e6�y�w��ø��'OF�+�^��b?
�K�I9}}�I���=��/H�w���a�Af�"A���JlWzcB�1�D5�|�0m���(c�gc��
�]��.̟�����Sc�ĳJ���F�)tE��5����|m_�z�k�.Ձ�#{.�zVVZ}����2)Z�M:��؆�'��|)/��[sdRY���9H�U�h��uX��\�B�(�s֫=r^�@�Hs���0����_��α5퍤->��/4��){���s��c���x��C��Z�#4����Z��'��)�*��sd4�]� M �ǋ��X?"��'5p��.�������.�[$퇒ILw��X��U���Z�\�\W���0^�J�_<"�D�fr3ƾ,�̢�����]����� �{ᅬjӣ������������11)~�)���v[d�S@��|�pXj,������V�6��Ufwth��C�N���N�����U98(#���a���6^6t%��c�&
��$wvv�&/�i��>8��ЛkJ��&{�f  ���n������Ǭ�h�����ކF��Y	�Rf0e5�^���J=�����Hk�ng\r������my�M�'����B_"���B���J�⇗/Q�i�p�Z,�FC����Ds� M�U�C��0��$�������VW?��R7��W����Ӄ����M;c� �%��i�5�m��ݞ������p������a����Ԇ�����@�y#~<n;��񀌡��b�R?���M��I��8ŸS�l�J�cP�]ӓ��(k����[ɹ���^�@}�~��L�<2��.�%v[��ac�+���s�ݺm��D]G�J7��ס��C�bMJ��^�2�	��������5�e�����d\�y���(=?$"�g�9Y9��TD����}<_���W��r�J3I�j�ݭ��A�'''W��i��{�T�UMi��*G�`��n�����4�Y������ik�	��._

���u@�������m��\~NMi�����d��<q��tq�f��A�jN��n�uJ�z����� ��O�����7N
Ƞ�Zs�x�~;WsI��yq�����>�)��r���������v%	�ր*	\����M���֞�Y�Q==��"}	��r�'3���J�nd�4}�jC��q��0<�f"�D�A���m\��rǿD��� 99vv2)g�H�rg�$�Ҷ>ał�`q��z�P�Y?�+(tO:-�⣭�&مď�y3I��d#�D�c-�^)������l+Ã��}�ωce��vn����]�o�����t�����n]T!��Ҹh�9��kg�~��6~V M~���N�[<���c�0�����h��e�����(u3�(��������������([�ͨfT���Ie�[������R�m���l����!��n �ԅZ��*�F��!��\ߢ�������g�a.E@CӤ�>S��xJ��Q��nk�5�"��]z*��QQ�wƶ���V����?ɸ�q�6��u��[�P��8} Q<��Hգyx�;������j7F�Fe�#G� H�
�v�~"���J���Ξ��
�>�����f\5N�;�0�Q��V��W�{�A���Y�BY}�\��ˢ�����g�y�W�ä$c�NP��Dp���[�0�̏��ԋ%��"�
�7`��ϲa՛Z�Qsr2
9��p��P�A���;(�9�h7��[���~�n�Z�1�]���^av�_P���X��/�6T��.4srw�\�;B�3'�3@���y`��- U{z���ڭ�뎁PI�y�)����\P��c��3��RJ��J�g�^$!�D�ؓ�iugD>~���dT$*Ǥ�+�5���=���b<�qnrtTz�Fߺo-6cg�����10A�R�U\"5 �k
>�/���p�����$�M��\{�p�am����P!���/�xoo�}̷T���
�5`$�L����7��C�w�2D�ls��)��Vq#�!!�>
���_jY�{/K�ڙ*6΅	߰z���<�j��61x�Z�㌧֍�ي�Sb��޾��V��d�TԄ���֩M�b�������\��h�.|uǺ�L�κ}u&{�y�����[Ǵ�`C'��PG��c2���2Vӟ��$�ס��}�P��lǙ�q�u�E�c�zn2V����ܱc���IvʁMB�E=>>>�
���:.��q#�a�gM�=֪=�����o�B&t0]Gj��^��0��*�U������/0������!�lSB0D���$�!�
�	��CV/K�U>��r��ZL�st�Io�Q���C��ds@DE���N4���|D�1�5��߆��`���
5۴�<�����k�M-A��Q��A��a��:%E�֮;� Fǹ#�z_<�TrZ�w����e#�>�����l�㲓���7Q(j�zg;����(��7��C�X�	���1�����Nv#�n���7�rF���^��"مn��h��B!�r)�\?���������\�Ʒ[�^C���m]7L�,�Gd������� x����8v�C�9\�k�����	����ǐ�Z����9�碷v��q�l�֣u� �y��Um3�)��b 0��-U�U�4�G���p��ZV�@$�H��� f��Oy�|[�X؃�.=��}�m:������.0{l�.�˥������c���d�36�:�1�-]R���b�Je�`�z܌�`k6��7N�)��^�э�������Oh��� i�:c�Z5: �k�4N[�)�W`0*"c��L��˗*\�4ow`�k�)+�����s���}zB��I����	w�y��|^N��7R��o��,k� ��U�tqq�a2	�Vh\�p������}������m�D|}����R��.^�0��n.nn���v��u��i?S^�8�G<����w�R'�_`:s��a~~����?`eE�<��UD�"�" ��OP|�����69vv͉.�aQ:�蛘\���F�ȃ�2K�S�����%jLd������C�0���s�r&�@f[:+`�w�f�=��;7��9m(��|Tʨ8c�W�x�~.�4�s�[� 7�~���>���?|Bt*.�8�U��' ���/7�
�㕠��7J̋�ኚ��A80̥�	�:�②,��4�[Xs��<3�~7���>W��B� ͝;�t��88-����+�p\�e#�g�B��Aki�F��㘃=s�7�QbQ	i������Dͱ�y�[ֳ�8�At���KF�K�Ҳ�=r$[���M���~��k<�F��1*q�2��c�n��ݳ uԙ�[��w�:�`g�I[Gg�'��%X�(�O��W�i���M-ޝ� �Xt�W��K�����WP]܄�c@x �#qפ<�����]W�p�Q���cF!@���5�.| @"Q�T.ϘY].-��X�'�,q���1�5�T�]�anF�;��_�f��Q�Qz&)�w&n����&��kzl��[�8��w෕3M������3���06�ç��f�K�b�B�B���P|�N���Rƅ��۝
`��v������ �=�	��:��j|c��߃.,^e�OP|����Y�&��M�S�!�.��H�B� ��>sB�ݎ�(m�?}c�%D�M��B/?K�5�}B�(2+΅�;�|j`�~x�qqٝ���u��!�f@��e�/���þp�;@�g0�-���4��/�[\�#4��x)�XѨ�؀�~�|�q)bz���ʹJ~����Sx�u�-ҟ�Y0]u��KK��\{y!Hbb茰����Ў̡�!�I��n(���#���B����'��`�:J�ŚW��}�0���9���#Gv�%��s�?A	/<$������qvsS��&�r��o�f`�T=�L�?s��0�1x�b��~�Z`%�������hJ�K)��v��5]����u?��(@��.?�,ݽ���!P,�Δ\Ђ�7��@'2��SÇz
����	T�� �~�����[�\��k��'���X,�?Q�"Y�L8�7 �p���Vp�LD3��f��>9<�9�;��4W��#�L)�Qƕ��1�j��-�k���4s��#���L�2�����֌"*c#
�q#�$X�Qy��q�0;
��55�M\�,��q�����M��L�������;{5�D1����ʨ�	���H$�!�TNO��X�2�����oYZ`YJ��E�k���qS,Q�x�tB��=...�bX�vZ�)�%	Bo-hƑ��ҫ]^t�gU��k��\�/���A���HT��\��\qu�Z���a>�J��I�.p牡X�ҕ�ݔ��o9�RYyq�ѷ�k�H@�_&A�+H�$�eV
-,r�;�"�i0Op����� .�����s,K� :�f;�E�<��II�PNٕ��I��WĆc!@kڒ}.��=^�8��y<�x��Q]�\�E��dŏ>[�/n$_�;���b���K�z��z���Gd=d�_3�&�
�eR�>�@������`�ް'��?���B�Ƭ�2�X�����ፆ>ˌ�����յj��u��kԧ�

�¨4��q��	��^���p$�r��<���~�J�!���r��IT�ރ���OF;�ŸЌ�b�*������Nˤ��d.I+��c���U/��f�3�2s	�ڨ�Ь���"�8ϛ����{��@~M�֩+r`� 3BQjFR�Ad+�0����2��`�?R�=�-���V� "X,777:����GT�7�x���h�,�p�ϕ|�quA/K�P�.�Ԣ���QQ:�_���K�&]�|��n�W����=X���$�1�ƘC��Ы�F�p�y�� �.��E��9fm����B����yfI�b�U0,Z$�=_OT,S�10�,�p} �_=gUE48�Mx�~�Pnn6\V_<ѫ3����P�v�p���G�C��!!F��S8�@/�CȰ��-�NT��zL���1�`fON���$������XA��_8d������u	���y��f�9�]#S��v���_e�!ͼ���0��N�8u y��w�j��CѸ��r>�D|�E%&�}zFy&]A��Ȳt���K�ܸ�`x��K_��2p�jlKKH�s7��ǻ���^9[���cm(└�aP:��C��E�.��Z[�����������j�����&�P�o��t:'�ꤨ,�RT
5!kG!Ր4��![�]�%ˉP�J��,�ݠ��11֡���`01��~����_�N�>��<�}_�u]�������ۗ�((8�δw,4=�.��=��$�\|y{g�e����a�O���0c{�%�x�,F�Ըs$��E���R�l��W�Q����r��������O-��|�����zi��\�ḟϟZ�{A�˵J�.���ik������s���@E�n@gS�t�`t�@!X� ����Ǜ�C�y��⪗[�)�feC�-S�j܏홥.}=5�D�rd�:�͛����_7�;R�)���%u��Ⱦ�~����pW����R�"�<sl�`{:�M�����WV<O7 r+�vt;�̨p�|r{AW���V~��SSץe���־P=>,���ޞ�5<-���-OR](�f6-���۷����	�R_�1{�X��7��_nJ5^�>�Ӯ���J��<�3�+������<#�evzl7��@W�69�G���70p:F������e����Z��h�����1����rr�룭ee'�O���SPg�ٯ��

f����������w��XwQWA����|�FK�6�%=���B�F9�Q���{�[�,#�Y]�o@ա ��=~���D�/>���V�����]R"�����$�v�;,~�|�Xh��3t���6��i�'A�fG�g�K������sↂ٪<I�%QI��Q���V<�����Cm�4�\t�� �[��i���R�tH MW�WB���5�C�j��.|ln֌m�.r���8jh$^����ء���ľ}�RS>����S�G�e�L&�������)
�*X�'��w��f��)Hצ���j�������4N�c9�[��xI�!4���b��,L;��u�ķ+�/�?z�YN�۳����pp���VffG�u�Msc[�t1GG��%e=�����a�U�p�&�m�̭Z��õȘP)�:���9))	��?�,[����(�R-���fJ7.q�r��9ʸ��vv����m���1�����^[���Zt}�����pެ
eؚl+(�SW_�~8[�O~�������v�e������Z�~[qu��އ����K3�ns��?�u��b(���Ņ1���hsf雛��,f�v0����g!�j�"�k���###���ή�.��t����IMYy�C�_}s�����a:���	K������ݾ��a�_�md�#ި��Yd�Ht���8��_9���Y�y4m�T�~�&��J��x����(����w�;$�������=���[B�ޟ6����騘��`��zT}��61.�W�CrHV8q.׽��ͷ�\���=�`�-i��9X�dޢ2�A�|!��(A�R���Ɓ��Wx5p���npf�N�pi�:1��?�z��4�[;<�YO���E��Ix��xD`���S�p��kGr��|�2|�x�Kk��77��n�*���5����NjN��P�/�	�<�4&������u_�^��.6��w�[YXD���wvG75e߽���K��^S`ЕV��a_�����z�����l���@ʰ���6-]*<�@�-�y����� �>�6��|�H�R��iK˘��8��	(�2���٬�q5�[�'--���"s*��|���e�Q���[;?_�����G�~�C����P�Z��yʱOK?'c�Ύ�e��4�طhƔ��o���R��Pz�c�$��Q�W�� bup�a���2�C�5Y�)r.���崲��
boedd<c�=�5���7�v�Z�А:&,�Mv,���~HRrr����Ǐ���-NmF���h�[�Q�=���r����Cb`���!�)���4��@�q������RY�
�M�n�%8h�n|�eB��sϘ\�����p�.�f|2�tjV������m/Y)�>��g_������cr���K��_O^{�89��oK3�M��܌��6�t{����T�E�����X��|in8�l-�"k������D�zW�3���
7�#!w�،gg�ڶm۬���{u%kQ���R��y�����Z	�?�lYDӂZ��Eg��H�����^����|]6�hhd��=��T��\_U��Ko�Z[�����w��e֣tg�,��|ƹ4�|�e۞"�����ߠ�V�雖�qȉM� �0�:�N$PW8 ��h�L,��ޕ�{�Ïa��:0�f�!R���Ac���Xܥ�
ڭqNDЇE�gV��F�@�ViQ�W	���0���t5.tuN?�JN��@�XC��Y���^׎��2,]������V3�����d��'IrǏo70�� ���[M�R8�����l��ƺ<L�-�WU��P��)��			��+6s��D�IL�%����;�E�=(&��N���>���dCqS/s�����J�?c��sP����֣T:;������������hY���Ϫ����0���Z1ˢ"##o@�y�єS�{rt˖-��L�SU�]^��8���XUmWvJ$q�Hsw��w����2,�Ѕ3�_�t�a�yF�7��7pc�r}���l�zuXfff�
D{zzt���_8�X\�rNw����Q�|=S�z�� �d�d)>R���5���֜V�����k�S���ựE�J�<��*O`��cTaٳ�P�x%�V<�9?�s�+�[B��P��c�j��$�ÞL�8����2:5�B�l��V��k��Uה:KO��?dv�����`�[	^���E��;37�M|���g��[��p/Ǡ�6�������+պ_��2�s�#��e�G@�rG��a�.�AQz�;�A�,c�˩��=J�o[���=Z�һ�t�@�inn��X�RQ^��0s�<�Pl.-���
�D��ϗ��G^^�ܒ�B�
��7|�S.Ek����ˢ����������I&�)�^��aw�SL�Qi	)��C�Wܥ������j.�	��#��
��a�{��ֲ�5n�w���=5���^ӟr�'ME�\�"8}AJ�Q��=E�gr.Ͼ���7�{Esz�L�˾�	�~�1��|���|�C�A�N���ȗ���zs7O\7fT��MO_f�A��sK�烊�V�����Oɖ<Z>H)��TMQ�H�25L���p�L�� ������ĪP�+~s�`ƫ+�g^vwuE�R�lk��R*�� ��B��w*A�����$�5���.�>��� �v��s���e9i)K�`�ҍR�08k�2�������-�3����TmV)+�B/0�, �Ɖ� ����rn��l�0�Eƪ�I&��!���/��N}?�O�9�L���V�4���)a�2*T��*�Lf�����C>��kв���]̡Ξ�)�㣇ɉħ�q�'M�iqd��xƩ��L�j�Rǧy�������.?��fm�*�F�W��p�,�~Y��,#�J]_�\nt4��֒rPjh]�2��΢l&���1xi�f%�(h��w�GHY�T�>�x����2x�\ӂ�2f����n�5���ӟ�j�/.yr���T"IoY%��T��\lU���k�rD�a�N瞺Ky[����Њ����2G�S��p��[@V���cJ�-�B�-{K܃����"�A��}�`��՗`�"������9��p����|�����ԪR߾��O��b~wѽ2�g�ީϕ�+�y��uW�*rN���jf���ܣf��@7�|h�2�:�m��Յ�*��Xڂ�k���,��#�RO�H<��*�k���9_:F�O�3��)�s*����=kI���*(آ���أx�����W	A�QI>�����L��osCc�즞=ل���3�VG�7��I#�=��;�TD�2���!ђv�����XC����/�L�s �a����\���(����s�jn�w������@b��`]$sr���I�#���6�/<�COZ��X��z�������e��B[�;�@�2G�=K�2�[��K�SaÚ� �~J%���a�c�lq���C���ma) w��5���<��p(3�e����=v@k�"�Ƈ����82$Z�h��	m��e���-[Z�1��L]�H$Yؿ[�(����˟kn2����j\�A�����c���LA�F��m/���'��Ř]����D��s�'m4���z7X3���a���[AnچZNY󷵎�C���y��Է3_
������-b^�=YM����y�:{�!_��b���ӜRN�mW\Y������f`8G���2g�e���=	0����9%�)�O��LHS�T.����fw�ݐ����m����q��-� �GOY�,�ฟ��HV_6�b��N撓���e�Db���@�<v?�����{��i @>"1H�XD���qֱ�̭������C�f���e�\)0�K2���_�4$�I�W�xE��ѹ�)�֛B�ۘ �M�����nT3�͸�����2�K��?����-G4��b�`�SNqUK*w)�v�dh�ق�T���6��C�u����*`#X�DhEn��E5��O���aҞ9kP�Tql���bs!V�v��L��f_�	ij�0�|��d�j����* ��N�����6u� Z�^�U
�ۜ�rg��ԡ�%�'�	�8�Gų�����&���.` K����H.���TR*9�[p��MLMá3�b��R�u��@���$~��N֧�ݽ��a��o;��]4s ����zCS���qw���<���v��_N3c%@_뾸�,�OD��b��<d�%|�Z�):T�v�p��<�߼\��B��>7����j�CP��{��� "q��Gԡ�������O�×b ��_G��Hj禞h<r�b��5W��7jj�3)� YasT�n'���[ ��T�$�7�H�J�`o)[N����2(=:�C��T �o�t�|�_vhµ�m��r�zL�_�It�����2YdL���kC\#&�l��9�lOm�*L����^ ��dr��@�6��nr�I]�a#��TJ�\̣���M�l���kn��v��}�O`?�n4�.Z�C�|�i���+���>th��� =���[���mFSa��m��b�ZEg\������"�*���� �F*�ڷo�$�t���ڛ|��7�d��������<"'7ݩvwQS9/��i�&H���7o>CH3�K笡s�|���Oc�\��ي�x�߈�n��SZ^�G��On;�I$��B�e��{`�}u@��+k����֣z�ia���-_�0�����D��8Gr0,�e�,NB�ի仱�z�1�:�?:::PrZ�*�҇o���;xh5 �Q,)K�c��y$�K��y��α����H �|���;i��=�֎8�<�u�\�>~7��r�:@a��Ī�Lt)<�+�x���~� -<E��� �R������byH�f�}��Y�|�C��I�xQ��Y�J���4�+�,i$����S
K���S�W��oa�⊣�j(�&#騸=���O+�6z�2�wbJJ$�!Ã�:`�� �H`۾�-����хpD	����1+�4�M�N���2O����u��g�`v!�.��).��ۚ,�>�>�`��򱱱�|7�V�$#K Gndr$Q���s7��b�r��x��i]*�Je7]I��E�x�w�I}�Wz�r:15�#)�M]�������13wF��p`=Г��3�i�R2J�1S�¿�Bר����3���B�u����y�o�P5'L⫂"��m���]�,��@]���0����چQȭ��m&�v���!U�!I�f��`%1ϛ�� �E,�wמ�c��WeK7�\{:vba��v �yq;{ج���?�li��c9�u'� ��7B�c�I=���Y�dO��������z��\s���I�Oʻ��?Z�K��(74����k��T�Qn>�}�Br�aXL6C�����|
&�3��s��;3��u�}2P���q":=��v�Q^V��KKK}���,g�H~>�Wu}b{�v�Um
zڷ�	= ���~łf�녮}ŉ�Q�[;L����Id�ʞ&�9?rNe��ɮ��zG ત$�)8�F.�K��R�LAO����3��h�ݦ���#ebH`�����"����8z��K��:���z�G{V&a��	XCG���3ؑ��Z�.�.�4˱�è+��0��M��������v..j���ٓ/K�MU�}S5�[1_���+�W�#����%K�C;OD֘�#���m��0P��]���!��a�D�m��;�`�ı^8�T�¼,B�}=��T䕖����S;�r����

_����\�F�x�� �Db��-�h��ύ�&�/�{*��O'w��+�Qp�+��ܽkT'�!t6�57߆a�?�n�	zMM����)+<��s%��zx���{�0d�=���Ѹ�M�!QM:�+H�Z�����H�=B�l�ɧ���C1��Q3��*�>;Zjll�C��~��JA3�$�U�B�E��o�儭�#Z����x>_��aAg��+��5�<��c###K��T6�
iа�U�b���#����_}���s�OvO��)���>����)��Q��xC����B�PŹ��ԎLIS ���y�>���i��D	�P��/����t���Z�2b u.�mx+���Yl��ɰ����9��C�o{��.��
I��j��kj���<�Z�WQx2%\,�cm��h́���Ka]�jʽ��� 6}A���0�O�ݠ���UZ��[�B��=ox����vQd���� �W"P��h3�9@�%=�T�#����0C>���Ta�|�d��^j�M}�r���Y�9�899a��Ә��F�1�X
��`�,��,08j�e���PV*n	E�5;kh^��� ��U"�j�权�i�f�!;�)����d!TH_P3���<o[D ��r�-�F�FTH6泲��f�� �~�x�)d9h���9i���M-նe�ݓ�0c�9%�C[�b��~z<�9�3$��G����+��J�*��{XB����"<�hg����7��p�֜��yR�2"�,�� �u� |�`��y����j���g$�%LF�����3��T�RUZBf�U���l@^�����?�^2w���$tK]������T��5�������(Rهr��S���f��$�J|s�^�jtv '
º�x=�I���"�Vh���|~llj:�t[���X,�6=V�Óo8)�^8zKN��s�$u*��1�xE�:$�G}�A�nBЏy�ׯ_o6ʵ�ʗ����#������̊1��caX�"K���̈�4���n�=vl�}Kjtfff�A�I֞bW���X4��c�[#r7 \C�V\�,A��XZ�,��Lj��
Z덠��ĭ��{���8:2���y�b&�8�r��_ϣ�t�� C��ya��Q����6|�y�Z��h�ژ�J�j�E�@X!Ơ�<&�~��VӜ|*Vc����V�^� �Q�YN�·cV&O^�P��~�s���IY4�?[؊��h_��v|�'ߍ�,:-�m�oIݐ8ӴY?:�20 ���fC�7��ֆo��+e�`��ڮ'+y)M����T�
����/n�S�x�x��	u�s�E7��+�o�)sH���!�����9tfu~�C�����$x�fc����jV|�ba��M���5����I7��9�4�� s:I���C�S�rH�N�ޖ��o߾��"K}E�\^�>Q$t�v��f���b�(�~-���;]}A+e���0��KE��*r�:��y/�]}J���R�2��6k(����������L���R���v������dȰ���w��[�l��z���R�.E��)���o6,���a9,��7��B$@���S�uN�eW�5Fqq[Щ��W����� #�\�<����^��ȅ_�Nf�*�z&����8j߬�ډO�*Bf )}c���˧T���`�4����XaKٱe�"���J�����8�R���oR������;�p�	��)�mԕ�L|͗����M��������n�p1���-F��s�[w=���([x�5�O'F">>~�s&��B�2���5��F����GPS��AW|��C�&[�Ғ��1�� ��QdmAA:�U35��4�`�Mi�v!�`�m�t:=̙����B�oN�W���A6��5P2��W��7��ʨ�8�J)	�7��qO48I�?T�6�Ec�hcc����G4��XDh�UB'�h+�3��ERw%FW�?# :p��e��
l���VM��;dGd���i\���"�����BM�!��<�ui�4�s5���H茀'p3���j@;��$�_44��y<L���cͻ�I�<ͫ��]zْ� �D:ج��n���P�����<#�V�L��y�V���q��?ʓ��v���]Ͳ x;x��bL:O�4�=��Q��crr�3tS�n߮E��$h�Tx�q��?���ؒ(>�	�HRH/o2�c~��@v�T�4oA���H\'���^	��!�]H����CbKx��4x�si� �N� & ���W��6� Fwz�����ox!�&F�!�BO;�8��: mU��7Qh=Fʖ��H&#�����P�Ԍt������1�W���V�$���|��s(YX���ί"cf*��5t/h7:x���E䅈�16�.#�S���A-̙^J�>���Lf9%�=Üa袣��>�45Q*�(:�g/QW��0q _��M(P[`�1�����
7�hr'�Zy1ncq�}���N�u�OCCZ@�� '9����^�ɕR�Ţ���5��+S�'�ƁS-�4��ҭ�b��9���IJ�7_Ns ��_����.�Bi׉e̡�)֪���f�y�&���^�L�@(�̃�e#[��P�fr��	��"y b�k�f�_��eY����嘬��
�Z�4N%�������M�����m��vq�CZ�7z�,��I ԠS��Lt�-f'qH�*�ů%ڕ��~���UC;��G;�z���9�rj@�rf_8�= �f�G���A�Xc�<𨁽��ކɛ�/l֋��ފ�f�?��&gp�ig+�\9P:1hah�5;�=��a�#"kdFŇ<u6���J���&S�SBvb����/�XRv$%�,��ma����5@O��������\4̥��Kۙ�T3h��9]]o��E!o�d�-���"J�W����8����s��nʽǏK0�@#/��S(mIc��)�=M�7<��;��M���>��mz��P��?JI�RZ=�����h�H�N%7~=e���J]�UR��ۮ�V|Sq�3�T -C]�_s/��`�����o~K��ޮ�d��F�2y��b�*_ϛ@TNp��T|g���t��>0�a��ѶPK4F����O�@�%P˩�u��ϼ�Yӳ��~j��fP�~#h�5O)�A�T���n����i��}�YUt\\,��S��U-6D^���Q�8�9l�'�zQ�����h��0����l�/�a���|��R!�E:w�k�I�$���p���K��ߨ�	^�[����"�^t�O��nQ�:�B�A�!��+A:��)�Q�a��&;Í}���%��Qp�����&�B��;w_Z�0p#�7h���1���[$P?zb�$�X��k��5��e�sO�˥�2�`wQ_;O0������GS(�a<�t=ЍX�ޖ�b��c`e�)
<2�c�s�}�����Хu���o�ai�2Yq3��n�T�k���x_9��ߑ��]�Yn
� ܔtceF��w�=���M�͵��HZ��1�_��"]�V��KA��"P��,�^u����T����p.�*��$�S��St߽O2���K(�| ����u�@�I�����r�ѫS���HA�V��~zQ���C�Gmm�������^}�x-�8'��\�A{���z��۠�pG^���K�7�>|�l|����q�X�k�pE���*7w��5��&���d)�7�P�P��*�P1�M|����Fݘ��XR��j�z��9x�L��H�m�͈��sH�E�֠�"?5A.�r���̲�O^����04����c�S=E�x/p�D"t��vO���)�^�x��?��!څ�����wM$) K�q���ec&�����!��E^5;�����ҫ����?�t��B�o�������]�x�)2%��/64 ���3e|�	���A�����z1ϛ�GC�����##.=��G�����/b\{y�,?�`�\�,ggϰ���@����՗24׶��~K�s3���c�-��Ik�=XU����JMЬ3�B뻌���8��P�v�-w��<��]	�Ç)�Og�^8$�.�t�-�Q(*.��G��-����L�R�(NC���Z{{}9=I�����A;v�D����������s�J�/_�~�����h�J8��)?� ���������@��X'�W{������]��H]��`*�`�w;g���ƌ�/꿬����I��m�蔾������ݻ���-BL-p������X;5u�իW�����6u��F�Tȁ��pHe���
��D�B4��j�p����P�H瞲��ȪJ7���%��_�-/-�$�3E��"�* ̹��\geŶ�2S	t;���`l��7Ͻs�s�:Q5�q��-@��K��X�bYK���9vnmoo m?+˹�9�K�ڍ��bK�� V��s2V!1yD&�c�>�k]�N��5�x���ɬX�R^1�Z�F�������Zu�Q:3�	���^�~��T�nW!ڐ
�\���'�G6˹	��+�Zs3jg~�����[����+�͘܅�n<g61�6ta	��$����ccو�����.SB�p�!����:�ؐG ����h�L�S�W�����ܻwr+�30қ�lش3g��Q�o��H���B�~�7��hȏ@g��gdr�uO����h�kE�Q�+&t/���##�%~l�a�-X��e�*��6 ϰi3�Νhra�N����Wхc�>%wz�3�{�-�D`��jM�A�D��!�=�GBSD�%ٻI
�5��#����U�%��ڧ�*��]��#� I��� �%��Ӽ֧�A&i������Wβ���Y�>6�8�T�wuإ�s��?�l����>�D���ߛ�9��׎<a�Q��M�_����p;����۽��?;�(⢏�,ge�rTC�d�2�� ��*��꛷�p���sO/{~?���?"|��X4z3�ہ�
����m>3����?_�ϊ�yV��ܝ
.W����ꔃ)���:K���!e��Ȱ�Txw��^8̏ѹ�H�� &�<��c��D�B��I�J����Q@@��H)w�������X�EC��Œow��P��!�RjJ98[�n�Δ���П;�a���s�8~�:]��f�I�"�8�NH��ҝvr���BX^���� ֣����
�C�������j�E�tg~�G;ٞ62㐸$�������6H�v#]�82�)#�5Ac����Չꛎ���zE#���`4�"��(�`~��{I3��L�����~�ey.�{������-��7�m�\rڄ<).�G{Z�M�t#�k2�O�������eLUnWK�R]i�����MU�$ü��v��BS�ΝIݝ�S�᷿ߕstu�SpQ	&s2�]�^��s]z2�x�9sje�A��=���Mr�M�IB��M������
�.|�r�K}`+�S	=c��b^{�\����>|J�8tW$�GsP���Fv��z؍�]>�6�ٱ�ŧy1p�S3���K\�'.	�L��+GZ�ǣ�omTA���@�u+4͆�k�?�4Ìv	Y��j�/6 %���-#��|���J�}��V#l��R"����wd��[�{z�tzΔJ�b���
��{+H���c�9������^'�\��ܾ��QϤ,7�aC�]2w�N�';��/>B�Z�E�h_�N�w`Wa��NN+R��������E�'~ExSY���D8�� ���V���3�6ю�I)\�2��UA��?i{����	�m���6�^`��o��In�n��Qx���uQ�:��D����F�k��Đ�נ媓(tSe�'P���t��y/3��ր&@�(�;�_>��/�rrr"֗|��رa�����W�̋��{�tKWBRR�c�O���{n���9����V��PwO�U��;7�;�r^me�����ߏk�/�<��`����$�#|x�tc�u|<g���N��d�MJ�AȞ�	@-GN�����)� �pa�2t�_�^��"��'�,C��r�c��r���P���1UN)����u�^���\]�b?��("��]�hq4�B1���V��)�|V/p1��7�qP��Ι(~/��3��G��&�!frYJ5gn
d�;�6$��#�--U&$G�T���ff�f��K�B�EEF�U�l��~Kkt^�z��"��a�ֳ�i��Җ�4c%�Y.|���3ߧ(����Q�/}2��F;��:�\��
7z)��q�v]���?f���ţm���q��X\?������t��'�Vm��5l79�R��e���M��|z�&z��)��+����>S3/�1�Y�?&��R����gc�����,/X'ly�����f�#`yϮ[v�&��Fi��X�f@>B=��u;"��I�CP�I&s'0*��Qo�:ۙ����:2���^B��@*\��q���O�+���pn�F�W��
q�_��閗���**&f�U��Q����z�ZJ39�K�Ts�\`N�xȹ����b'���I�����LL�@ЪƓ�����2~���H���ZVU�BȎ3x��Hj���p���<C}3�X�E���ˢ��<cI+�K��D��6������i�;���ߚH�Q��ke�u����O8
*xX���	��cޅEEOu3�D�[G@նB3���޾�i�0�6d���
��+UyP�@u�D����'K"�N�O���U�i��	.7@IE�V����O�f�|��Q������!c.��5�1h�Es����$1v���Hl�e${�F�Yvq곲,T��d^*��vU)=镏�o�N�%�V	L�d2��# ��W����Q�τ� �i�>~�W:�����3�1�Q"�2W}���h.��Q:����ë?�%KiM��u/[����-[�Eƞ+�"E0�*W����B%��3Ϯ�KoIN���g(��t����?x���t�N\H$�m�Y8�Zdg5��q�\�^6=�_����XwL�C%Oǜ�s�rsp�Y�b?�8d	=QZx0���)���j8��/�~q�Ι���͢p���(�#k����W�*�Pt��v)��0>��Z�^�r,Bn��=(��=�_Rx����&��_1q
Ӊ	��T7Z��aip*q�t$���rv�0�砂}>�lX�����?.Y-.�H����z�'�B�	���Urhׯ��i�t�A�l�`Gw�?�꯶��I���V��'C*~я�Ȩ����?�qk�>�c���ۓ���l�5�D����������H�j���-��S�5�Y|�|�)�1�/�ʸ���o$���!��l�J�Y�_��M:WEW3���58yV4�X�q��������@4��3`O�`�׀P������� �
:12�-��5�:ѕ����)K]�;�k��!7_�ۤ-��k�˗uLx��U��u�^�;��ļ���d�)9v�=~�0�i��/_2퍝��M���g#x��(��4tc��f�u�F񈴽mD�v�gm�[Q��}��7���`�s�5(�LG89�?5��U��N������acɢ��k�[2]�i��PU�|G؆2"k?�,s\\��/���j)�Y��B���9����P�#U8����G���J7h���#��1 1�n�Ю�H%�Ĥ���!���ѡ7�dj�<p��J�Z;�s�qo��tb���i��_Me�/���e�ݔ�D��������+�h�Q"��T�i"I�IY^��_Ey�:3`��xD���T`NpU�ڑ9�[���̘虱�)T"�#a��k}�[b%�2<���{���`hVX��?|	��-�kO�&S�{�;S���~Vԍ�QMh�BT�̠8�X�g�G7��vVcmFj,i8 L�3p�	{�x~fpvq/n�ߤ�Z�z@HH��K�{���#3� ͏��k�{N�bA��S:mxbq�An1ɻ��)�αTV�.}�xU�*�l;��^�{�	�Z�ݱ�H�|䖛Q��Z��*���;��y�LJ�a|p�X�cEs��L�i�9�Q�֓�>�֚�}F�wtgH�[�!&ּ:s[�s+�_A����n�O	����Pȭ�d�����~��ʅ�OG�;�L��A�ڙ�`���_j|o^T\|Q�6�a��W�H���o�2����ATO!��5rg�)1�/?L��ib���z��k-�9��Kh>�	��&��Q��w���P��#���Yo���W�������RVl����Vh�X-�4���q�+ב��A��N/g-�mpz�5>]9r�>�F��i�M6PSxI����a��y��DED~�E2�s�a��Nc=�~�		<RWٲR3R%>���d���\�MD+ʾ�u2��$j暛�knް+x�%?Y�!1�����6;�q��c���w�T�gDl"
:��9KNMg�+4p.B<ƑiM���ͥ2w��UL��?Q8t#�_����*����6���!�����U�u����z�Դ�y�pAI��ݝb1s��Y{#W�4*�	�zjiXƏ�� l���)��e��az�˯��*8;��$m}XA�0�����*2)�!-�$.eF��q���L-|���wo�h�Y���%��A����&��\�]��í���t>1_���_^�ˍLL�������Pfo���/!&ځ&���D�����(1*��f���ڕЂK�x�U��G��3�q��o�	Pu02�ӗ�B���G����DFOs3s,,342�h���\�P�q;v{t��ه�j����]~HNh�+������^��G��`0��E��G*)��绰8�k�j�o����vI������qP�'�����䐩&D�e���37��By�L��@��ԙB�B{ky�����]��0�"qkB��[/3X�]�-T1����m�**���?�)B�m�l ⫟Q@no'�:��y^���rv�(Y���"���h�o���05�r<A|$ݨ�T����4������2���Y�mA�\z{��D�Aߏ��d���ޮ}����R��n�7U@C��� p��Z<��GF[5'3���k9@���L�R��Wa�������5g�N�����u�۪�6��gƚ�
FNW�&C��|[||l�V���L�np�G.y�V*�d _��Hx�g[ak�p:C��UNь�;!��/vrқ�_ p��8��`%T=�{u.xI�7�͕�͠CSf�V(�*�
�I��;��@~5)�V��ΌWg�Ţ�;"�;6�1�P}����P�3�o�}�^6I�1 �,��p�T�m�޼��Ј��� ψ���͔s{+9
u?Pl��L��8k��&.D���z3Q�w�3���j�3��N���64�scn�������j�Uq@v�U"c.-n�FX����+���}k}$�+�q`�\]�ſ��q��)ux�dT���}�D&�x*��+�w��^"{�����"���$�y1���)�e��|,�5C��l� ��_�{Ї==Y��x[ۈՇ)���z��|���#0F��٨6<P�ۗa��J�-`6�ҭc$BbH�YC�9��VV��o�wc�x,�,������O�9N�G.��m�꜇��G�ޫ|��� ~�� ��]�~�����7���k��������Ti�s�b�E��	��g�����H|h��IM��j��+��#�mޠ^���&��sb��+V��$"�R�uw}�O��X��+wwu�{��+��ۥ�H�~��.�]ۏZ���99�ҍ��s'�t�:�XR�|Bn�H�?(�f{{�����aJ4X��\�m�Y����Y�T�򾧟�֔j@�
é�Y�u®ً�ń������Qr~�����	n��Dl8s
�ܔ�EF���X%�f$����͹W�ޣu �촥Д �r,�P��!���^SKsprhs���9�JV�	���E��/�w��|��o�>�����	ݼ��§͋W�8�$��k>���!�]DJkw����z�a�۫�˦�M>h�?B$��6S8�	�TyV��G	��ߗ*�����J��o�`�zD�5��@���zb(�+φ=�}������G][�T�{�uM��N�@!{�F�׍a��99�����z_�^�g�rή���qx��K;ِ?z��emܥ�yU`hha$891�;�7T������"u�b�Sл4��mV��@/�%tE�[��]Z;B(��^�����_Gw�Ә��������e<��.U?ې[�靀2�ҳ��$m��,��p�o@��q\g,�U�q����l��,�e�]���ЃR���ǯ��?8c�$�Tq�_yU|6b��K���4"&�S<d��s']��9I��{a�mxA��u(��t�3�IVu�Wb�/Mm8c �dw6���/[��A�o�\����1i8$vZ	���T�r�[��j�,h�|Y!ˏ��Mꄡŷ(�N��L6�J��/�T���s*G�Q;@0 @Kj��o%��x@�Yz�	�����}-lu�]b�Ui�[��Gaq�w�H����љ�%�lH8ʶ�OrPJ�p��x	�6�|�:�4��8�!��zkڧJIq�:�r��'TT�q����f�a0��ݏ��8۫{u�lv�2��i/Oz,=�������T���Ф{|�%�z� �j���nVk�cն_��~&�ދ����l��W�[ �)���4�1��V��6��Y��)�k�r���3��-"��|R_����aa~,�7)�	�Ώ��m�I��#��v��I.p�ĉ�]�S@��kmZ!��?g��ӹ���^F��,����]��uRJ*&��(?K/i\�3H�#��M�u�_�EK�ZG�p�HÞ��Ƭ�Lf��s���B8��_x�NH(lSpo��0���o��be�!������Ew��֛fi�O><�\�J(�㶷�z��.��+��8�!Cdu�.��&��ۮ�G%�=�m>6+}4�B��.��R{�C��
�:�$G�/8�dw���&���~a��^���]���\�ȝ�j[�7��Y�O\��@�/f?���lk��m��}�3y1m4�SH�X�Ԡ�ڮ ����MQ�����+.��3��:�A�I�[�W��>�󭤆~���3T]G��Y/\��]�w��^s:����iOq��Ch���^���w��O�4�S:��x�k�~l�?�
T�'4
�>�|�Y��7-�!��q��\�8ipN����Us�m�c&��ܺ ccc�!!zt�;S��na6��-N�7���3(�U��>g�jao��1>�����r!�fuɟ..�U^=�k�/�s����|���G\6�?����W��ЇuC�#R��G|�-	��S.�/�*��Sl,\���1\�d���"&O��>�F>����[�5���ĕ������==���$�;�4�7}K�k�^�P�NP�)�b���$~�n�͐C��}Ƞnۓ��o m��|��jϭ��#k��gf��XK�г���|稤5Xy���'��kg��6�9�E|��*�#�:}�(5���U�YG��W3��+��nޚ�˝�!p���1z��
#��jj" a���S�f$O�̩����$�Z��&B?ޖL�>��6�Ρ1��<��k>�J���E�2h�p�@�1��� ��'���mU.�e�Y�A��ۛ*���J7��$@m���DCcm��>K[]\�q-��p)� Mv��B#�0VCY��j���S�Q��5�lIrv�H�K7�ןݾ�G*'�-~㙣H���\���z�:>�f�Gn,*[-�����z�K�YR�j>U���y0��t̷+Lp���?6o��ٮ�uUQ�܎���MiG�!�1u��ſ%��Vt|�x/��6��ݕ[��,XGE<李EO�E����/���_T�S�'[��������?��b��j��i����꼫]���WK��,�z�tds�O���ѥ%J�y��lՐ��9�I�<�R<��\WG/�8�z������Yͥ��&�EUà]��^'F�����T4��6i`�@�y��NO��w��.�{dš��>���&/�����"
�����o^�cX���;���&6����\IA��q�O}�%�CW��<��O�i�-��t���͐���2��B����;����7��VPGA��ڈ`T�`1"��A�����Ju�t+̈!��!E�AJ$JҤ�B��|?����u��de�˓g�g��>{�s��O�r8C]]ʮ�bRB�깡��ῒxju}	Q�y�v��b8f�������g�����Bj'�'`�ď�4*o�J�z�Y� ��k>����\���w�i�VVT�}m�_�Կ��������N���H���zK��dݘq�?������̄=~^���O&R�@Җ�	�Z���4��5*�m?d��`!�)��<xw����A�Zn9�Wk�rKl\N��ݵ�%s��T�U� �ݒ7O�'�x�Q(R��!~	��6[q��R���~������ ��q��m@�F%b�C��"�>y�x�n�ҫ�tl2��ϙ�� FN���i���,~T��U��e������ߞz����Q�8��E|Ɖ:x8�" �h��:�I4����X�UV?���b��ҡ��X����g�r�������g�M�i"6��6�a��7�G�S>�>Žc�P�w�ι��r�+�/���pE�����C�����+��8شc%�Ĥ�Aȋ��f�M ��S�+_��^�2���KQˇ�"�yp�j��Ɍ�d�({E�ZˇF���-)��C�r~Or���]v��
�+l���FVq�&��\�/�8R�;�Ԍ�p��rB�"�=�_�խ�)KWX���B�N寅t���W ��Rp~�5�(~v�ο�4�X/~�Yu1qI�'�F2��$cd@��)Z�^0h'_e��ysGҖ+�ޢWazf���q�����++��F_,N��#In8�&��}O7H��J��#��=*�ͯ����Љ�2d�������$��~��NP�DR�k/9y������[,&���$+9�K�d�xV���aYWU���7?vA���։��|�`������m��Q�J��(�%�n���Uv�Ck�i���1u��Q&�w��>�(�Y�ē=22��,�y��zE����@�az�
ӗ֌_*�N�#/+��1����=A�?�������)�F�  }�yW`5�����7c����ٸ)�p����X���������ū����7 8���,�����7ъVnٹimSp��*Bȍ��۱�G��J�g�d4w�f��f���(ﴃ��"��@ 9{[���8y��f�/v��tCQG��B���j�Ҋi�	�:�
M��ϰ�q�ħ.�Q��,��e�{��
�J��u?�L{`��-(��*�1)��ҧ\��$+�� �J��Z�5Oe�*5 �)��p�
�.�8{҈�!X�J���8��b�%���P(^��?/�]h!EC���H�UͿ��T���]�@�d����t��?��7�8��BFX�z��)����m\r��� �dL���I0w7����A�HUA�eV4u^-���!��`�Bk� ����U:6.�m ��K B�d�mB���,&�-��A�9^��;���o�1?6����
k��:��_Y(It�!K�&��@�p���d��uÃф��Θ!e��H�	�G��ς�ZQsk�����%�C��N�˻�:$ѳ����
��w��F� �� @�F�R�<N�cF������Q}�,
<��w�@�$��SE��
H�F̃n?����ߚ7�0lp���c���-	��f��,�R���/A>״��������6�����0-�M
<���]��T<L��e}��s��4����俗�� ���a0굍q����u�e����)�+��/�� ��R� �+^��U�����ߥ��
��}_���(`8��e�`� A��t{�P�����f���!"�d$�z��#P�]EV��%�9H�EUz�pӁI3h4Ȓ�f�$jf􏏏?�J�A�b�Q�F�9�uG�\��.��"��H~�։# E���ws,�-����u���w~�	,�����1���l�-埥�}si�-�m�������0�-���A�h�%�P���h��;Y��#5�֣,��\��	`!��~��G!E_>K��O:� ��ew�nGW<�'"�t��Hdu�D�p2o ��F����]�.�� >(I2(��dl��j��Au�wVՈ^�Q�m ��������ʎ�:CZ�,�ͥ���\w�3����� ����9�@/�ZrabtDjU;���8G �{��$¼�4�;w$Q��0�K�oP{>!�!k������	���Q�M_o%Q�뭴�n�+nuY�@���-���Af�VEE�n� �TE"(,N����J��f�UR��;|e��!��bEÚܵ&�$�e���D�~4 ��dF��`��&jNd��1MT�6��:�!g�e�M�Z�f䡽ԅ�~��Wf�s�%KV�^��]��ݘ���+��9�_����ƹ�Y[�;Eod�d�-��e���q!=�	��ȷ���:/|�l����Q�`���D�MV����3��W�#�fe��D�g��S�h�`�N<F26}�yz����G)��dD��[9I�U}��%%%`є�H>�#`߆�VF �2x��൲ׯC�Z���yvDYE��"b���Z1��y3*��]T��n�Jj���qR����ZW��*�b�˪u��M��s�ٷ��6P��F���WA�Zn��1�7+Q��G�Y|���B��iI���Ew8�G<�.>T||n��g�?�>������J���y����H�Y?�˺��i:q5��k5�#ȆF�ז���}_������9�\�!!�0�k����Ю�HO6���g+{خ��F[���猪�#�������{�u��K��������QUo0�A�R��ؑݻw{��@t[��N���s��3�֡��w��2��2Լ\u����p\RtY��[W��F�M� ���nj1�ܔ��w�Fg�v�Ai�~�֚�#��h�)pzF��D��Y�t{�+��k/�j$}�%(Iw�[�~&qX�{�Jl:`�]IlW�ߞ�����@��̈�.?ᅗ��<&�#������>9ɮ!6	K���pT�)@�Ź)�����@��޺×���ȵ9���d�-�qj>ӄ�ϐ̬A ZK�����g��@��?��O�#N��3��neHt����}�K���׏B���$P<ӧ�{����,Ev�m�3a_�}���z��v���98{�w+���Ht���Zc��F�S��P�(@��0jT?Y��x�$M�����I)8��0�H�آ��Z���ĥ��>�X�Q~���ē U|�<��:��G�O����>A�������}�A�}���5��3�^��-�w�<]�bʜ��RZ/+�I���=�/�jż�V�*z$�v�G9��f@Q/]E�!�_9T�:1�[��=�U�g���-�3�M���ǟ�Aj}��G�����>$���?��,e,�L�� s)����$yb$��Z۴'�������"�J+�,w/�lb˩4h<�����4�3?�����A`�Q� ���*���9�\|"����\ 	!����Q�ɸ%op�M�>�X�]�ԛ)ZZ>���6�V�ҩ��[;��1��	�gAY`�h)���ڥ&0�ϣTY����܊
ڲ���]�O?׳�cIgh��s��>�vfa��,��c��yg��"I8��>['��T�~��T�.
�T��8�I��͇e�E��u z�Y��ݐ�ġ�m���|'�
�kbd�A�tz���$X;���_��@�:���;���ӸUrx���"2�:��O>���# y]��{�
�f��\�}DMf|�&~���z,`���u9�����<j:!�5��K���9 �X$�����⑕���?������}�|z�j���\ZÈ�6�$H���g�P�qv���'^N�K�~"A��(�ϑke.;|�����C�#�������d�Ê�! ��.�����~�W�]�d��	:{�[Q_��Z���b��+U�Ϟ.6��.c�
Q��7ܬ�>r�jއ��ˉL}�g��,�7�p��*�ɀ#�[8�xH��}IFyon��M޴+�zk廍w���ξ���_�,J�BK %���섾�`�q���lɆS��YXu^�I�kL��'vd_e�1���GC��Qr&��@���o���̓�a��$&P��L���0���LNN������}V��5c����/��ڋ%�2��6���G��Րj�.x�G�c/�ս�8��0��_��8"񘌚�x��k��6QD�z�qR�����Ꚛ���oQ+�a�:[��40��6��a�>�u}i�}��`�(�\q+1I}8 #��j�NuA^��ێ���݇�?�]w�Դ���֧����Iޟ۸�d;$�2�%?n��Ã�@����;�ۻ�W�f\8�&���k�&T�1@�j�D��c���k�$�O�8�'������	C �H]#���ߍċP���D&��� [gk��m�ȈNa!ǝ�T+����h���^�٢�F���\)_�zw��:O � �jx���<�niI��OL\Zٟk#g��:E@��Ja*$�s���H��2'@�	m�-����%�Di�c.DV�y��L��f,²���X�f2��0����K�Ǐ���2�������ك�+/�?Ǧ�3��*�-H�1�,�-X�(oB��1���0v����u���`��j����kpDxxڅ�Ja��N�W��|.^�s�U��ԙ�I��dm�Z`[�����ط��U��"ӻ���']UrU�ML8��n��7ͧ�����]0��?�V�WGf��g��͝�ԒY�ل�!�����b ��D��L�K���!�n~�C�}�8�l�8�gΎ#d��ޅ# M()+�����˫}���r*nu��p�U ��z��g��Y�Y����Ӌ�)bEe�":�
uk�=$�=�Hd3~��W� ��4��P��GN�ED�NW��7�ǩ�U<	�������#���u�;�Gq�j���l8�^��n���4a�7�;�~k9I���F�h6u�pp�i]��u�y�39lƄ{�H���nؗ��"���ܟ����`�1D~��G��#q�HksI�}]��3PAX�C�ѡ굆4�ӟ1.�)�W���<�i��NN职:�*M�����3��+��.ɍ�9�w/<���S��6�U��"�����u@;}�	/�������	p&��{����]���2���[��G����bP�G���2�{[�����/3����?��ӃhSki�ㅬ�[��ܼ���>�Wk���V�?D:V�u��s���ݸ�� �V��5.�a�q�j����'�p*NL�dG`�9��0D�s#�u׌k��^�_l��Pd��UL�ƛ33a��ᣥ���3���{{��Ig��&/�zEi��]�7k����"�1õl�f7{��O#r<T�rz��ʕ�����0�z*ֶ�*�'�-BM���u�q}�����ټ�0�@�-)�LV|�a����	L�X�s����oe����4[��s����Aov�S#M{b��c����v)���:��0̞y��[\wM�$�5!\���<�QK�b *�2�%�3f��¶�f�z������bj`]�%�E�\$�n�����#�R��n1��� Ѯ���mq��9#��z �<R���V�a"�\�;_�ߔ�-	!]�j��!��ԫ�}���{��'L5��?�1���Ev��VF^8�^�2��+�\a�	C7�ٗl�cT��\Yk���6?B	�2cц|nf��["�
�u�!�c����c��M�%h���OR0����2�hJn���]sA*�﮹QT9����J�.�rF����o��B�7�n��VDTe��Yԕ�]3	\���	+���CSʠS�����g�p�Z`�k.�&�c&����>��D�s�R�ʹ�U���\x�!|J�Yr���{��"�s]3T[��{W��G��;Iv�n�-�Z0���BVe,�ZA�g��K儚��!L��U��'���l"U�Q�`�$7 /k��m��:\�Q�a\_	c��[�2��,���
��{~sl'	�NĪ|�n�$��"R���R�YفT96y�1��L��c\�O^�f`�a�{t'Zź���w�W=�B�������0"Ùb��W)����NDF:�&�Y9�{j&�8���:��j3i��O��g�h�W��:��R�Y-��T�e�
�j�Y_�5yY6�z�j�����<����h�F��Gp�uj�pMÏ�����ܑ�D�� ��hka�B�l&��b��]L����V���Ϥ`+3{G��]��-{yxhTd
Er����"\\�[��b�z&x�Ӏ��%� �d����׌���6�������P,o��Bp�7����n�ָͤ=i����X�Ǽ��1~(zt�(�SƈL��B��:��6��[�g#Xmq���DI�T��Iʈ^%�Y�}l�cH
 �񳙰�����g;�J�L�-�^"�����Ԏ]ų�=�T\G��wAQe��!O!8�
�S`��������ͷO(W�M0��Rnogg�p��t 6�'$�8w�=6� M 8�ʁ:j�ʪ44����(]F������Ʊy8�q��f�<I�-jD�&Q����俟4iT�|��~���������X*�D��W���N=&�T8��čj����Ij��$�I.�\&�Lr��2�e��$��/�.�C N�f��_&�Lr��2�e��WI
ٍ�N���;�qC�Fn���7��8�j*´��ҏ���T�?�~���������#���	.\&�Lp���gs�%S?�V!���I��<��Ҏ��Do�C�?�]r�r���'�k�Z��&�~4F�+��ѫ=��:��BM�L��4ū�P����$�0�Q��7K�:أ�-��#y����/>_�����rI�:�����j��Uc���e��UI�?U,����;�(��Q�=���÷셛=��D#,l�|a~��� PK   �x�X䏆ze� r& /   images/46a4a336-cec8-4b03-9de3-7f7682b07e1b.pngD{P\Ѳ�0�0xpH'�{ �����kH��������!��ß�����USs�{��^�VqN����  �>KK�  �{  
��>�}�T'imW �l�����W��7I-7UG7Ocs���'��������9���eƉ 1 @	�,!��y���ef����QP�8V�&�сi��j�dЅi|�`FI�^Τ�����퍘�PKXl����Omّ�؍�^��Ѱr���x���n�f#����\��Y]G�\��5p�HvE�h�n9߭w��w�w����6E(E�~�&��bzXж��sh���($o��qX�OI�\`#������;�uR�.�is.�˖�����Zt�v�W*��k�E,yh�c4�O�g�AbИ����{�{*�ix�^�������� �x3����v6�k��w�jZ��-���a�e�LU����j�������
n��t���E�^�!� ���W�Sul�emd�ώ�b"�b����E1z�)����
�\K�F��2URS�K�v��؅٫�E�E�;��7�|� �ؠ�cDC�gΏAT�&(�J����,-�2�oc�b\��H� �C'*֭�Zʄ$���H���o��Z��z�QXi��r(a{��,�_�[��R�ˍ��جb�|$�Ȇ(��NV��(���d|��n��Ik�G�?���(ċ��	�dHpG��Y�OM���?y<%�e��X�PNa\�vs�����oc��������h��9c8�=8��PU�F�cbl�>(&��A{o���1<� �Rhg~S�h{ѡx�GCCa��\p�N�R:=_6f�1��iE�ܾ5.̢��ِ��Ve22�4{�U���L2�Biv�k��LCM]^'����dQ� iZ'6�e�夋�'K�����-8@՛�S��3��0�2�z�f ��K1�
��.�}Y�F�7G�O��ic |j���0+
�q��+�B�@��1-$��q���Y�R������젆�]�]�S�:S�N�B�����MSXb�[�Y���/�
���<\��	Շ�ڭA�pS��L��Շ�����A�>�p�1ht��"("�Kx ��va[��R�t�R���
&�L.��:�^8��#�_��v7�����p%2ơ��@6�������Jy��&�]��+ ����·- -o=��F�DML�\KW7��b�=�b��p��Y�\+��-������
�o�DI�k��t�R�LX����3c�T�3��w 7b���NB��/o0�� ��t��ͨ��� �fB��Cb;?��S�7A-5\y^y+��~�]g�w��/	��EQk�g�q��R� �fm�M�Hh��F!��f-����n�G��H�>�k�$px��a�j�ޟOX�0sx1%2g�p)i.ʤ���xa��Q��u�؝ ܲ�"
p�zM�N{0ȥ�{����\����P��ި6KR��A?�N���/jc6s ����u-�b���rH��Ծ.D8F���.��_Cx�GʂpfG)��8j�Op����������tY���O��+�ޖ�iJvpM��A5zZ�y�������"��7�tn��m�O�kR�/1DG����0�Ϡ^�E�g�x�W��M��^��w�<E����3$su��?n�PZ�v�_�3K���v�R)D����Q$+f�E��P��5��;���@s�y~K���@WȂ��x	��=�"�c14�X���⿒�%�ffef]���	�����K��Nm"�:�R���j�.�
�C��0rߪܮ�����/��*4D��eRy����'�x�/�89QQ��jx^v8O��T�b�Q}y�T��QZS����c��Y���$�x�j�`=���h��@U���"���B��f�*U�V^�9 z>D�s��:�ZL쌩��3��
�_�9-|h,�ޙ�����VY%���lm葼����?���s�N8��Է[�gXv��V>F���Y:���TL㓜�ggO�6u*�DY�I����^��*�1����Z�T��|4J{�~�cQ����F �pF��П^�����V�9�k��+@��T,�ԃ�j�S�o"��13�Ԥ�@_Y��Z$�$�>6�͟2�87P��0hWP�Gi�:G�ړ��\�Q`nX��`�`��9��*Af�/�� �%-2�8���WA{]h�BaXfV;?j&�[--�����g��n�A�C_&0���BQL�#NӞy�]���AФfLV��V:>BW�7b �s!\eU%'�Ҡ�?�[�]>���>������n(`�[�7	e�:0a����d�ɨ�^����ܨ�I_k��8X��7���{�Q��gEY��8"� !��\a��|�<�9������9��	b�JjҒ�x�b�� %��7��z��^�'�_���[�dZFF�Ȅ�a����"�EJrr��*��t�H�ßW�!���79-�n�#��5.���Y�ܪ�5�t�y�0�&,{�O҄S��=�j��بH��Ǜ	?��-�E����̳UE��r��,D���g��1�J�q�O12{�/�u�t%p�f32q��?�.����A��;���	��A�I���>>C�a���+��
W؊�[ϳcxa����o��Ν�YM!��G�0�������4�e���Ѭ�|G�����1ے[P���J�F�ǲަ�UE]3S��(��Zgw����֐6�/G#칊�JχV�2�+��>�S1J�}*�`޻6�Y����= ��V �~;���K�GPTc���H5�n����;6Wq����Z�F��0��_X� �8�s�cG6���Z� ����EY�F=pH<�S��r�:��JW񛃪E���yo?�4����{>�ͧ-�gk9��a�+��F���]�����HAD�9c<���ܖ�:�.G�:I���?>�O��і�v���3�p�ϰ�ɼ��n:��۸d�`j��^��T��8z-f��V��s�Q�b>X �y%]�(B�@���H8pWw?�v�}�Dds�:�CؒXl7���Ѿ��a��[�x��󂐁��*.����VA�� '�7d�|u�Wo?�v6)���O'�q1�;�؜����W��=�5�@z=X�}-V91�V��>J�z��2�p��O	�1`�Q��N�I����t���ڱeH�"S�Fm���)|5�[v;�=(	���=����T�(�3hXUTo����G��u��S5�م��#�/+�pB�< �����8���L�Xw�[�݉��_��s����O���EӓҀ�N.���r�g�g�D��{��F�[�T��A��?wӪ���!����iS�-T/�Q؃��ˇ#
�D�*�+�>�6n���ڏ���}���́�n��bOھ@��m�_[!iCV1Y����-➑����N�����0B��L����=�79i��%�_�R�5@���=���"��݊�H��TGN�~S<Y�9F�g�PǥMJZB=�d��"�H�ćC͑�p�|����eP�\��[P�(5��>=�C��9+��W뛟O�qO[��:- Q�{vq�8V������N,��G㎯7�9,)tDA\k�S�}2X��^�q�l����S�'۫}���O[��ݭ8x)�
�BW	�� 
�}�Ȓ�V\�w��Z�F�tK8>� )܅����EI�Ռ��+���)X ���*���&�]�\���y�\���V'��KF3֭���#0x�k�3S~��
�5�Ǩ�nLL[�H����`�ŊT�
E5,�f[Kt�(ny:C�OJw�`�����_�J�l����OhϠ(���=�c�t����Q=7�/K�!Y���5�o�h���T:�T�����U�)�7(\�SS�X�:3�|'��=1�g
�v�_	���@v>��*c��<N\q�cc��J�ɪ�������pąat�T?+�5)��5QN�Wbt}
��>=7
O;�_�k��68����\�팕J�9��`�x:�<y0�|���P��xV��r�0	5�0`Q��.���X]�������R�Ws_N^vt��Y=�5�ۭ���Ʒ�1�Kę�c��4m?7d$Kٱ� 5��X��*[����{��[L�G���IKe�CD�L���S�ԏ�;�I,@B.��'�=����f�wC�Y<��q�e����������*M�%�_���≳/Ӑ�a,�q��v{�胬��!�jk{oY�A~f�w`k�4�~}�@�k��93��N�����p�D6#�Ce�Q��U������X-�yܦ�;}�y��Ӱ��݋-n���uB��(�C.�ݏ=<!"�P�cv��e�<��lct~pһ�*%�Ǽ�F��Et����k�I��E��S�R��tC��,�#$�����VJ�f��W��_��o��̀X����!�����8�R��*��*A�u�j�A~��{�3&���$���˂��V��
�`"J���C_���ȱu��=���#�뙰�#2�i�A�����-��SW.�;�X�[rc`h�fW�Ae@.�dJ���:�w~�R�߳���]T|� �u��Yn'Y��ēܯ�uX�L!��c���Ӿ���G�4�1����I��b��IwB|`��J�Bܽ��p���O�`��Hz�B�$ϻ�T	QVY��6s�td��%�	�<��ڜ�ǫ9�M5V����ZU���?��Ƽ�	yJ3��o������r�Ŝ ٽ9��n�:����w��g�W\�7����\��ܟ=�Lߠ������yX�;1�r�}̏E�W^����d�y��}��$3��F����%tNB��|i%(�wXP����Gړ7~�̀����﵍�iLө��^zݏ3��1�{�hϱ�#پ��A,��2���g�Mo]�I^���7�RB�����0�z�,�"%�$�+T
�&�P�63���8E�_81����" poz7��f?vY���䛎�������4, ���v�ռ[�82���� �8w��.���_��ٞ��&%u��Jޢ� נ ]5��G-|ş��ͷ�E]'�������!��UK�c�#�?f�2�tX��ͼ],���O���G�T��H�#��P�$*�r�����ǧ�x�g��d��$�d�Q�?���7�-���,�	_9ƈK�Ru:�mG������0���3]��N;7W�U�r߮�;�&���	>��7AQ̂���c[��`�C� ����g+�^3��p~.XXC�?(ށ'u���@��X��j�&�QH	><i{p�ga:�r��}�@�Kd0�����4���dh�og���	s�-5��9l!u8��[#ъ���Xa�&��Դ��{v"����TY�N���?{�\zo�5z<����F7��0Ꭽ+7[Ƌ���%*H�/�Pٟ�}����jp�� w]���\�{9��P�WuO�VWKt!UBj!'�����jyCd���f��V#��Ρ,~]��ѕ�������ˮH, K��=t�D��\PFMj ���h����w�"�j��'E�Di�؜�+}ӷ�y�|�XX���S��u1�14���T\[����2��pZ����E�dY-��|{���u�H���7<{�0;ʁ6 7]�}ԍ'�ܤ��[�����S|ٸҦϡGp�a;��+h��3u��v�T8E*���99���!>�X�kgû\e��_W�i-�������V��Uw�#�g]��w�%�J��c�a���ڽ�40�d�-)���d|��X�b!Q?Z%�}o�_�'٥3VɧTJE8����-�]�ʄ9_�z��P��:rh-i;�{K�ѩ��S���r=@�ֹ�舊�~�ܘcu!�̝��3���&�ml5�m@��ޓU��a~�y�~5�,/A�4���AC���H�6����)���8�w���XY���b�M���U6�j�н�+���KE-��N
P^�VT))	5��`s�Dt���R�Y��`�ĘC����>4sO1$��E�o<�v��j5�c~9�E%�e��c���#��2=C4�k>�{�����8���7�>�WN��ԯI�J�0����H�H�S��1���n�?�j��rMT-pRhG�t1Å@�J!{B���yK �
�ʳ�&,Ü���o<���ؚF܊:F�<N�Z���\��;"�6�z�ړ=ˈE*C�4�����o�y�������@;��bQ��|ɖ3O�b~_��Agʢ���Z���Ag���vKv	�끤��¤��F@�:���C�7}�e5����'�ؙ�,�c_{&���d��"�6O���ʴ�������՗K�E�{��L�4�����9���%�����7�����h�$�]���T��)�"��D݅I�WM�j�S�����^�/�X��H�2_Uz������ǭg��Ӻ��)�Y�5�t�(��ꂪ�����}AKU3K�+��<��F���:�#1QĽk=7NKT��H�[���9�_�9���O���乊�L�[	c��T�t�$f{����L]W�Ů�x\�ԾV�L�I�3�z�u�v��'� ����!ݔ��p#�x��O�)�\g��o��CY�����lz��u��,��:��f�٤�-G_�v��$I��/񯳳lu
Ԭ{�>�lJM+���ԩb/l����=����Es~jPW�A��(?��Vu�
-�hXK��\�L6�n�O-֞C���^�?v!V�I;w�FÖ=^$��Z���/z����b̒9�ҖO����B
={|V���L��Ӣ��&���F�&W\�	��et;��!Ҙj�ΐ��C�[5�C��c����b�ؕ:�e_�t�S|�5�R�t,<����i�ȁ4s����-��M.�����ͥG����xX>�%a��e8�=hX���9}��v���W�
��W����<{���{�y����q��b)N��k��\c3E��4�-;���%N4%q5��a�akjVVǙ��M1E��k��Вkҳ�Y.�%hb�-Rݏ: M��E��`�6vN��O�J���"N֌�������=7_����ջ�7�~CXO:+�D��ئG(ѹm��:~���@sq/P��8��Q�`'?�FH�Թ��z�_�c�i)�\�� �[������K0�$"X�1v�6xI��ˌ��3<--M�><��]��E�9����J���pѠ��I���  LŻ^�7�B\)`)A�ɣ���Б�a�9MM�8}�M/g���*v��Ң�^�:��M��-�X86��>DIP���0���¢����Ea�A�z���]h���'K�K��[��Sy/�ͤ5����v�bB`HN&�<3y��p���+]��S��:*r~�R�����n����K�GE\ͩX�d���W�	)�m�����g+���(M�#dh:����ox�8"1#x�;s2\I�乮�C�AhG]86,���-X=F4s�:�

ƥ��)�ޗ7i�)�H�<��[���rZjL�K�*���Y��c��o�JS��;F>ı��nmm�����0�mі�'I)�N����9D� 풲���8��n@j���g���&�k�FV`�9qi��ܱ��b���PĐ݅�e-wL����;��ooIt�Y�8Ͱ���r�E�C�N6'g��_�r���6��m㠭@���%�S��Q�-�ZN`�!@5��y݊�3@�g쵲��i����OT1qq�155��CS���������+�y���LH;;C�,}�[�Z���c�-e:���u��`@/B�l3S��~zh �$����2.���)�=�j��| Op�fª�K "A=�v|��B������C�G�ݡ�؆/���TQ>�y5�/������iXK�lp��A��RE�y|AUU�1��?m�#��Pg�jl߿����9���V�s��B-
Ђuu����}d����W�I���$�������_��PQ�ՙﾁ5�b|Z��x�ic��/�D��`~����u�#�2��t��>��,�>V@��_Z����_]q~�.��Ts��?���7d5�,�����yt8Li��^�D.T)c⽲g/����n���tiR�I����
��i��j�ϞE�Q��v (�USZ82"�!դ��Q�\�h0�� 4F@�t���_���t7��@��ɇ�\HM�/�،�5f�ؿԿ�);�����vAA�z�L��M�*���[Iʷ���וe�]W��}�39�ц�ӿY^�h������KJ��&g=����#L��R��oQv�V �'ӻi�X��_�!�ݫ
'��&o*������\2	��c����At y\�Ǜ?�_S��Њ�W,9AH�{{{�J;h��]�޼�����m�[~���u�lv�bH��%��GNЭKک��xD���d�Ɗ�����iKI0A�����ۋ��o��~3����{����tq���`��9d|0~s�L����j*�@N�Yᢖ���$�-1Y-�a%nl��F���ө:�+Y�w�.�D�U�Nb" ��T*S5��2��Μ�`�9�e� uH���ݾs�������8��oK���q�%����Q�c�_�d��$�@SSKGZ7Cŭ�6�q��Z�; ~�'�����(��H������fܢ&�w���_ �4���tϝ� ��k���y$���k��b�:�Li�7���P�>\�Z�|�x�c�X��dQI��%Pi)I������햭�x;"��̃}qB�~�m�PnS�GM#�<쇇�Oo�����;�,~�T{~Fiw:q��-nyA�}�O�4˦��.�%��,���C�G��o�`�`�^2�0~^ ����P��gnG�����	]����4�>&�0��Z�#�U	�o�Dlm||}Ơ�0zEde�����SB���B̤��'Ύ�Q�}t7��F	'�uUL�#sڸ��a�N��<������]T7o;�F|�]S�����73g�蝽�"Kn����rg��)Q�����c��` ��F���k#/�3ɏ�d��+�o19�&����cQ�/���Ja�:���@j��-���i�"GA�XZ����3O���a��J��i	��Պ�hf��	5ֆ�����y�	����v�]�DQ����p +Q,�\��aذ2�oqݍhlVE8K���������ֽ�,VB8+����zF��y�����o�u���!+�䶑�<,��}�[�u)�K�ò����d;UfU���Tzu�*�|v���V+�c_RTJ
��h�n�]L]������(��q�u�ie/�{����gf-�c6�!W�;Wiy�xB�i��Q|�K��
aqq��������>�)@f-xv�ڱd��ƴ���*�Ъ)�u��Wm	\�8�Ɵ]��r��)1���׳U���fG~�.1�XEO3��:4�c�q��?�F�5<̤c�k���p:�#�ST�(�������@Q�;l �U�úrm�3�P�����2�W��ZP���Rq��O	��v�eo}Q�*�x|����&B*�Ckmm���k:�Au\�ᶿm���19_Wk��-��sxtm� ��A�tA�}A� �����j��C��^�t��#s����k�$~@����ml�o�!�9�E���CM����2~z�����S��`W͏A9�������Z~;�j(��ύ�a\O�l:u@���]��c ���c�̰~�6gR���%���j��Pm���d���z��Q����ꖢ�9�����]�w2F9\�#�B��L��<����4�M7pnD�!�b뽅�F{���b��CqMM�X�Y@�� ��k�끇���6��,��M9W7�.Q�䶍��,B��������{��ڪMW_�]����|㰣³�7�� �Ĥ�\#���n����f�=`����?G���}gIk,�(�#�c�8�D)�F޵V��QNd�[�����*
���&�lG�]�N�guu��F����!�����M|>����j^��C�_��[����JUA���J;�\����"?��ˢ��l�}OY�P1�T :��W�_�k��	 �~_8.k��7��N(�`0��O�axëhs��a�#�GF(�jl��XW	�ྒྷ|�v�usX_��#	I���TO�v��P���H$��1�����f̵g P�%�["�n(�j���"mXW���Ĭ�˜�����{��L����A0Vѵ��,p���ņ���1��;�Y(+4@ƻ
&���KJJB"Nfg�K�8c	���)�cq�+ qt������X)�(���7]ٕ6t���k�+^�`j�=����qi�rX�w�N�L��輍�:K�TSƻ��u��G�L��yy	(=X\K����:k!�7x�2o�?��p�a50�0�k�G����v��A���hN&ش��	�vd��[�[ej
��x�������+������y���G�%��gܞ��?��m��N���7˗�쩖���4�����I��CE��Tjdķ��ȇ'`J�BY�Tu�zS|��%���6���l�������������N����}�|��-��v���Cr��~� 9�6��K��J&��-�T�ӡj��s�+oz��WOdV�M��'sz��˧<!�ő�7L�f&�����Q�Viз��F#e���׸4�D�:�}ʙ��:><"��06JY-���rwA�M �K��#���w���(]��u��t�Tf�֋��Z�N?�~_^Ttt����|��a/.kB��C�y�z5��^����1ܻgp�6��&%��s�����V�i-�_ɸ�LH
�w�Z�3��q��Z�?`�䀽u��FBB��ݥ�2E����&��?�}9����ΊI
25��=�2�a��ݯCwSe�����-��T_�/�-Gz��lm_���ۛ�;���I1X}��\H1O��=??ۖFb��v���S���>�C���G���'k��T�w\kϏ#Y'gd%$��Tzx���E�F7]](��ߒQ�'bՊ�YP��# :��ˏ��ҋ�!dg�sM�P�w*үi���6=&ڽHni��/��z��F�fl�R���#~�~z�Ʌo�4�&촚YLb 'V�g���^��t47���Mk����L9yĨ����St�^���=B{�j�ҩ(���7��W�ʛz��j�pgy����tG[C[·�5N<_�P(g�UB�fG�8�}���8���B�S�m $;�\���9'�6�Ykm����V��n{�l�:��K���1^��:f�����&�k�}�>�	h
��Iw3f�i�1��G�1������M��I�����Qگc
h^{�aL����qe�4"L�vtt��$�@���Y�9?�wP��U{�W�a����Y]]+K����<^j��A<���������ps�f��:O:ao �~�ar}�5.��{e+�Z�E�#����N�9�ށ�;�nQ�>ρ��y��w�eW`z[3�]%xu���^�+�����B#\�Y��&f�mcS��|֬����bԸ�\l�1b?9��{��|�釔��ꛎ:9��葲���]Ş�W�ߑ�b
0x2��fX���`��h��![�?��eO(����1R́������1S�0u�	`�t�<��ּj��!�<�pb�m�;Tm���R�����1*9��&����.5O��8f�~5L�c�vՏ�w5j
�SQ�T��}bm�v@�r�`����fo��߳�i'�oc��}���:n��������ֿ*�˼ñ�ս�Q�+٬�G=e�d�D8!I��� �]�,�>�����45;���x���%�� �� �7����pl����	�A��$�k�O������n�����n�V_�o6�a�y�������3�!і�p�A/%%5��8K�|�'"��fޤd������mA��P��
Gѝ�Ֆ�?91pn����o�݉�x��U�\�~|�y���&W���I�M�A��� ��xx�s9|�%ـa�Aט�i�JM�}2)&�-lV5�z^<>Y�]_]U6sz�@)n��N��XҴ#�{iv��/^t.t3�&�]	HUV�J3S�ƫ˄���:��.MĒ OO?�+�jEBᮏ������n�v��G��̲c�)�d�dy���=i�w�bF����=�j�d�L��u��b�s��<�ɒO�J�)�u;�pLw��tKà9� �kUj�'Dc-����h��o1E��f1��C��7o�����Ɯ����3��<bR20Xy����R��?4���w��~�����lTT͏�f9��a|薯�}�ݿ��	����cgH�/)M�8�	��
9f�s�f�pc<1���/����I�Gv�������k���e�ܹ+ d/����r�-�z��X�V��V�d���h��+L'�7��vL.Q�f���������]|y+nt_�aT�.f�$��/�Եk���b?��:������x+�o�cA��vZs<��ge��b��l�]Vg�hj�i��x�~����+�-iZ�:J�)��1	a0���d���2!�9����s-�"p��!��Ч��^�_Q#ȍa��)�����@�������f��0;��GC�����ӹo�Q{�m>����7x����~�PK�L�"��Vf��@q��k��#�qC=��?�?h��md�J��O�DP�������l��u���6�L�*5�Kaբ1wIБh���{g
�̨��<�sr��g����s�*ӄ�n|{�4hv��`�Ly�/mt>G?�W���S-���DEE�ޙ�5@��+�1z����5KhB[��1��&L�������ď��׻�n�ȗF:��ə���cG5d�U�@��>�\^Dd�GK�� ���㋩^=�Aϧ���C�e��GxI�$������F;Jɶ��H�Q���L�Y�^Ao��t �����pW?�s���P煺d+~w}C���O�[���K�k�z�Vq�2ʛ1+$>2X���I�K��V�n�
�f(?�Fj�R�'���Z+���=����Z�y��yc��S�"0:��6?�R�W���o$ ��@h��wKF}\��i�fө^	��Ke�0�c~LU3�?!�i�e-���Ր�������9P _&vpK2��!�3Ȍ� �_Wb�[�f]0\\���QeӪ�[���O0�RcF�|���i<��U1��wt�ܲ,e�̡�����e�����-���K�|�I�3�� �氠oܡ��K��_�)	����C>�+bd�/E��kN!"�V�A�!�6������]���&R�Q���s�Ͽ�k�t]�HF��<6��--��_�w,��Tr��J��a
V�[�m	$�B�`��!��J�,/��i�@01#
�Q��H���>�/�9+>E(�|�O�FXU��Y�,�B�M�5��ק�a�\��Y8_;�����@�����5殓���{���䒗!ɥ:�̼��A���"5HT+��횅1�]�~B}&X���j�VY3�e�JI����Y��Q�V�S��nd�b�ф��N�^���E�.���9��;{����e�|鵁=x�4 įOC~4�kmk[q�f��@"4�D�[yC��\�:�/�2��j��,�hkkz�i#3w-�~5�**�*B�9�CdǌnˬA�o�s#����wd ��Ur0���r�Wz��6�L��/8=1�'��L��M��Qba��ˏܫ,�x\����Cb7���z��2S@�#e�AN?�}Y%�sW�v�W"��tU����y^��uƔ��yZu��r�c<6�1�Q'�y,YZ��B�ׅ��P���[{G_���N3�J�=FE�|�0�_�>D"��,�A@g�V�Obt(�vt���<)�&,�;��w��H���,�ַ<��.�Z9��^/�&���A`����4!l�I����3Т��Ϸ���[@��[�eJ��uI6��?�lB�Z�
�9ED�����իKZ��F�X6j�XV�A��78��^�R�Q^װ�u����>���Ն[��A�K�S!=��eg�N<�p��CZ���E@0�&i��q�i���b"J����w��n�ꓯ3���#Y��YM�׶E�y u�����!�|�n�����?C�n��u��+&P�c�P���s��o��ͥ� "�0����٪�Z��/1�e�A�)a��~���lUA���� h��
Fqs�z���q�&��;LXCN%:!��
�RS��N��0?����Q�����gon/kM�m
�]E�z�f!�.�&�^���8;�Q��6�������.�^����`�2d�|�������d]�����e���9]Af��W��3�F�a�j�<5��w����դ��+�<�x�a�NmŽ�̚@K�>(9� F���X�������sbS
��[���f�3�+��j�0�0NkR��m*Bxj"���_2g��ѷ�?0$RchD<� o�-�=9h�:�u�-�(9���Uj�h�st�1$7�QP��3����65���L�����ma(�D'}c�l�jk��\
�����w� �S�ZX�������b�L������"��A��at�*��r1Z������4���V��]�?o�0o��8ѵI�O��jkWA�(�ςP�8:������0m��w�y�#]����������YVW�	��*��V`p��&DV�>�����s�:�&>3�"�O�r.�'^�8��I줪�"D����!��V�ׯ{!4J��g�ָ��k��-�[l�t�?��x|tN�%�'o�\
S���U���G���R�+�ҷ�\3�$�u'�@$@�Jjb)�~�.$��PK6b��x�v���1	ٕ7O�������=恿<8a�+�:9��O����K"���E���ב6|�WA�1jʌ���q�h���\�=���� %�>Bx"���������7~S��,X�
��xPC?L{il+`��]���D���<���f���M������Cc�l6�?i��$G�W�^�.����S����>e�ܕ����h�Yˀ����ߥZ|�X����㎻��Ⱛp��Xď��`�H��G�*)M������I�E%8h�,�wd�D�J卯��(O6�B�����,*���e@}�F���`�c��L�|tw[u47��p>����������|��L�m��y���3*��V4u��$x�壘�!A���I�I����n�[)U�yL����������#x��3 }��h�%���?��X��{��{<J���A��hK3���QE5�w*��4
Q�{�Z�t�!�V�I�}�4�e��=B�?��\_O<���=���/2x�e���e�@T���˳���Lٍ� Ǟ���:���&�0O��L��JVv�a�VU��K��n>�;��z��:?)�Yɉ9��ـ�{W�UK��gL��a��-`/�֘���HЉFT���$V��%�9�%�y�5�o?��t�����I��R���H7�󑒨��5o�8�}�����<�(��F�q�8̯�!qU��U��y�]}��cY��5Ɵ���|�y�7Vx���-h@kF�<:���#���P��Iʨ;Ƕ�OY�Z-��9}�ʤ�Ёk}3�Fh�_��N������xwN�P6]c�-d/$���O�>��);]�DdA[\&N�u���5��i2ѫZ\�f��/�����odZ��C5;n�B}n����.���_;Ĥ�}�ADI�"���VB��R������ZQ�s�(��_O �¸��؂ȶX+v�R�.�c�?����<4�Kѝb[:[�58}m�	�0��gN���7�������{��W��N����bg�Y;��\���Lh�*d:�������.�����#-L���j��ȴM`��fc0W�)?ᤡM��#��無�C��t����5M\qt1
]L�n����,�ҳ�e���<L߈!�����5�A�G��qo���{[�{|^�"\���H�f�;!^�7���x���&�Nsa�z��'�3���� X�δ����	3UJ8e�܏�?�����r"�Ą���Ξ�)~��b�$�W7�A*�.ن�'�k��L�G����D��e����W��j���҆{c�c�~ݲ4D�H�`9�OØ�N4���?w�-c��?���ڹ�k,�������J��R�������%t*��������ց� ��U�H�$��N��:�k�i�W�� [�k�ғ.m58,��ϰ��,�[�:�����%Zf��wS+F�Rh�,��g�3����*ן��"�&H��ǤR�ɇ]短4W�4�;،O�~��w)�$�+)��V?���X��vߖ�������p���A�sU�>����!�w�L�86?�G��Z
�~"�p]����P��M��6ӄ�	�N���ʊ��HV�$*O$���ͳ`�s���S�j��^b
89�w���%o�"1�a�^��$�؁�
�[�^��.
��������޷�"-�R�ݵ4�Kw�����) "ݽ��tI�Hòt�4,.����}=���3�>�u]�3 
pxhh�*4�/^��&9\�ց���~+��9+�g���l�K���ExS%<n��D3��N�=LʆnZn6��B�{-��kHڴ%�d���GEZ_<�_=����������iO����j����}q�����5��g���)�P��K�:�N�6P�/gk��$���.ઍ~tYN��I~s|&$��N<��d�Z�o#�2n�/g��\zƮ{A5_����a;�`�`h9�U��_�Y���_�@�;���g��+7C~����*C!��ʷ�ߣ�
�^�k����S|���%L�b�Qx0���ڹ��]c},9=�f�(�D�����Q>>��+����f\Щ�R�H���;��8gD�u�ZҮ;I��?=�����a_��l��� +�3��ۻ��B�/9����� �#����S�����7Ta���w�6�Ѡ}�6krә�~�.i��vr/�eѾb�}J��~� Mm���go�ꀆ��8l��j��~0�={1��bd�Z^Oo.-9��+��w�]OYk�w�3v�WS|�;|\��[rc��Bt|G���^|��"MiO�P;�����X�ͫߩ�������Җ�Ӌ�Ӣ
�������is�j��J��u� ��|yBH��$�u2�,A���:XX!�k�.1#,���O�U������GnRQ�W.jXRt�[��%	^s���<qݨ���L=���?�5�,p�vreJ�b(�^f���JF�ީ��3�@��ۊ����~̽�u�����17ql7���������V�A�w"���N���5jHb�gum��ϵIu�ʺ�$�iU�kF�"ś����4�l�C��<gZR\����3��-�lBO8hs'7��g����$��e#��	z
����^�k����]m��-c2��z�껴�ߋ*����@�w�\��5�^`k+\�k��yǺc��3tΠ�;�tb�r�ғh�x�-�cxC�+����x��>uj�TP RK���@��A5�N�G��±+�W+y�'2��v8�:oN^�%�z9|�"j���g��i�Yէ,4j�E�%�E��X�\+s��n�}3j����0K`�R���r�z7� �rn50�9�����g�������Y�m������?�0?��1B�����@��y���Wǂ����-W��;�iwxr�7޵�e��.��ooo�6Ȓ�C6���'����Q����Ny�tԃ�"�ν����LT3�`̬�py[���ЎP�MA�H򌞥����L�ǫ!����%��;�9�`������]2����3���猩�����qf=��g?�9uw?´���\޽�e�nLtI�icQ (����3�v�o�00��J��l�/�aJ�	Q��p�x��~�l���oֱ!v&
0B~��d�z��j�2(�߈�	�ᤲ17�U�U������]QZ���F����J�]v�B*<c��KT�c���x��!��0��Ȯ[x��x���L�h��#���Uj���p�}]	�i�C>�F�x���O?a�ׯjT�ɜ�0`f��o/�6�L?Q6�m�-����	1����.=�4"���q�0���A�����Vb�B1-!��n��V�׶ QΜ@��V�C��r䠉0{���T�|Hɱ�y��:-Cy0����xc�K�q��4��uRRRf?<ks<OZ�j��Ͽ}o��_.1"v^�����w�u� 8���I�@����]��9��iQ�lr4��d��ڟ�_"��2N,vn3���7��ǳl��x\��Z�����ܼ/a�#�Kc�~f��[	���34m�3���7���cޣ-�ϑU���}aVz9�'��/=tϞ��I�{<�����NEH���D3�ݮ�d������7���">��E�<��0k��s�Z��TӲם�aF�Z��
1Ɲ�S7e�??:ki`T���|�X��kyh�ޟG��[��p h�]x�����V%���R�@6����-�z�|�������b�pu�Pa�۝'�q���9nxh�;�-�eu-���;�˓ո%�e�aY�rjr܏����xl�G��L�+��I����ݣϺ{u�A���1!��3���������4��� nz+���e��9b�ٯ(�$_Q�[��
���cܫ��g� ��8���I}�����#u�~��}���v~�ZS�uDY�K��AM���9d)��x�H��M7�MUa�9����A��^�K�_� ��[F�9d�v)���J����B�D�"�>\dGϹ��CL��w�L4�:L�ʕ���e���+�)w�E�F�E6E��2���S�����8�L���G��K(na��s';��0��,�#��9++3'gIqkfw���y�����}�C��I�����)6:
I}4Vu�I����R��%b�=#N:?䙪-we��B~o����r�n-�p-9�{"ǵ/w ��r
;/C�x���A����_��Ԇ^�wL���ܱ?��8�d0E��X�y�ޠ)�ր��4���?����25��]y͝?
i�	$QS��P���Й&9�u�E�<=Ymk�\�Ė"Eŷ4��2;�2��� Z���J���reWM+OO�O�i�i���;�ѓ�-T��3���o���أF�� @�������dɱ��r��m?[|
�i~�%s�񙅰�K���n����������X���]�<�-i_�ptt�L\��LL�}�6�G�?8x��Y����Em�t�&宅ۅ0�6���Rg�=�>��Q�r~3#N�Ϧ�UI���R�h�H���d����ep|uWkXIDL�aj�ꨂ��Ҳٸ��� ���� �:�����YE�Fm��$ڋS�W~�-e�P�,__I/'!�g(�T�t6���01{�q��~`������fe����mI�H�����i���[m�lBPl,Tl�''�<��Y]�*��ZSL���{|K�����6�nK���<�ͺP��肻���'�(|�ɌV��B�A��fɩ!���<��n�cEk�D��NdK���	v���w��K<蔡��V��s�7.!���y���g��� G��x~I5?v~N��Ȱ�Ur��(�)D�n�&Ђ�t�u���3H�|�XWaY� 5:ra�������*b�
����#n滂���䢔x�q��*�htZ����*�����͕3�8�[}�&�D�����ȍ�����Ҳ����Y��S.��=�ӑ�g���٪�~�'y� hi���F%!�����o�C�g��{�%�8n��(�����H��W��D'&C�?U9�M�Ѓ�\�Ve���eB��g��d�������M1����o��
�=&�u{-����.�|T1�>G�^-�ga�oBp�����0�M�.�����_���
 �ubY���s-ak��t,�l���{8ű�$@���؏c޴㼅�����`���&Q�f��2�h�mm]�Z���me�������إ��ul�||_+��w�q�QbTT�=<&���7���q),,,B��2��'��A]�`*	�h^�1��2J��d���dA���NH��K�(i����cqm��!������F^P��Zp4���[�[l��0K�7БC�es��� �~M�(����ۊ9�v�YeeY�;���;A�ӿ���;����i�^ �踶��C�1@�#�i5�G��% �W^�U��}�sq[IV�%��Q�]��`^l�L�.m��\r<��\P?�Q4�B��]�! �r�σeZ��x�ld�,<,�Lٞ	^���U�X���l��zxz�p��[�%���X��r�9�{��+��؜�&�{���Bt�g�ܗ��&���1�^&����D��3�~G�yO�Q��|���;U&�ps��a���]�ON+Nm�>��ڔ����P��� �F|��jL/��)#d��2U�p]]���	�v)�I�?�M�2�6�7T�d�y��ׂ%�؁���7���;�7c]�Y#�����U��zU#��yǟ;�fŧad���\���-].yC�^�W�6�0�Yq~�뵑�q�U�w�&�x��;6��"'��|��EV*"|WfĶ'W��6{ueM` (�i��I���p�3�,^���[���¤��?6p}Ӡ��K�Qߩf��<S�2ƈM��2,ȇ�OJ �ĺ:�V��|���)�9�/3>^_�ʍkh�s%h��2��EN� �]S�
�)D��ւ�Nk�Z�Mp2�9�2�������B�[����'�����F.�	
����>�м���Lby&D���'(��L���<���)��aT�ʴ���:2���k�s�A�(2*
r:䦃�����������@��J��M���(倎fH_>:GQZC�-��_L�OYC�5===S�;;����do�foa�Ϻwttt���r�~���%��\�&(�XT��4��1�8��� \�q��LF�[���[\ն�e/��L#����lf:8��љ����`��bL���\�7z���(r��TL+�8��TL�g���c3J0}}��@5�'� >I����T��P�M��y����gjqr�~^�`b~��k��g�C'y���+�/7�������%M_*�lzi�(EVt^���FXx�t�(T����4�B#�.�Oz�t	�B�ZD���8��u�����Uk�d~Y�����mW��
�ٰ���tO� Z/;I-��l�I�O�`����� R�k�/�A�99Ŷ���n�*gB%���s����E�
�ccc���_�bE�DI,a���,j��%|wΈ�JK�u��DH��+���/���é���(/o���D��k4��4~���q��H`������u��#�n�"��SSV?��_|mAVV���
�l��33) �DX$�h�x%�ށ�x���ʕmX�E�yd8��Yդ���*i���d@ǀupF��$j�������	�o�;iY�Y�״���Lʛ�j�aE�@�W�h����V�I�b#��6��a��Y�F��ެ�����v��H:�X<�2����*�#����9xwm3������)�A�����}�����˛���A�^s^��J�&~Cǐt���� �pWZ��	��VD��72�2qrε���9�q����4�7]-j�V�g��؅)��j\7������N�NW�O�F���;���哫z�]ʕ��Ĺ���11¥�\�=]�����u#:�q��m�K�a�{�_CA������Q��e8b�3�}aL~A��������M��d�~�Mj-!�r��%%P�c�򝥯��APfi�X����5�ewf�b�JO@G�����o������̒�D�<3V�0��R"]�6B�T5��N��1ҥ�Zנ� �u�����Y�@�4򘕰ڢg�����5�ZN_�,�)qήrU�!��r��f�w=��G�<܏0׀?��	��1��4�>(l]d��Z�jbV�s?p�����c�w25Ӌ�q���P��7��Y�~��P6!�,B��+�+�q�!��"ه�Φ�~����
l)�����kOOx{�/�`� �8V��$���e#ះ�x>��U���L��Q���G��΂r��*�2�ii�b{{�.�Mo�Ļ�F���H-4�����"C:@@�_�Gͦ>����~�w8ߘ=@$
O�s>�wqq���������e�@q�E�@�����8Ms�>�@KôKTF[�����]ê��h��6h�1�'�w"z{��r�zr�� tˣ2H��@���ڧ��ڒ	R\��D�M��{H��	<��3���EsB�_����%�iL%�T���b�v�Lh!2��FR�Lf=�Z�`��j%�c�+����s{ Kmj��$��w�7ѦkE��Q�����;˧� :9S�^STZ^>�)9)����a�jx��z$�x&0�����6�g5�#��F�����xt��ࠀ�	�-�#�N�؞�|�y�Ӡ;�Q��
����-���`0g*��H+�i9`����()�\�&7#c��u���X��Ǿ��i�w�T��F�,7�����L���k�ޱ�K'�~v�K��2ZP���׎����^��Mә�Ȏ��>S���8�c��[?q�1�N:��M<*:�E�@4�>'�LY�S*������tH:�,�Gvu�9��?�d���K9k2u9_���q_� �v��_�^�nlUA�z�*?N��ͅD�������͠F3�(�L@�W�	��G#��P�R`�8�Ht�!8�v�����6unb:�;����غ���g���W-�pnLI�߽��@К��˲���}d���!��{��T���Vo����o;�HK:�ԟ����L�0j����7�Qg��VW������������u������4(p��ɴKJ��8��mi~>��+��t���1%/NV�_���uƘ3��G!6�Ǩ����{����ɸ�w��\a��"vT��;>���A�t��0E��$����	R�<cJ�}��U�(x
�h�-���^�=�G������w2$R�L����~�u�N�fݏY]�o��3��XӤoIt����H�V�xI�`rg���z�G*{��@��?�����Ks-�b��׃���=7�����v,�e�&ٰ�u�T�V[)�u᳍t��n9K���}�78!ᵡ���<hU���CSK+	Ć�Ļk��yY������[-�9ܯF�ݩ��2��'����`�����o�;��<E_#VM��F�L�N�(��ᑑҲ���:��\�rEG��I�Z2�\X)3���E��'Y/�j�E�(@����̜��������I$�����NZN���#*��]�Y�����9��\�L�Д��m�_\\�ď'��9I�p�?(	&$����{�)����w@d����N�5�s�l�h�Sj�H|�츜i��D_q��'SG��sm"_�l���X��T?2�Hb�ݕ�������&	y���&֜�ﾾ ��l����cq�WN�������G�]��\�Y�9�7�X��R�����4��Ӳ�r�9�!�̾D�}j��Hd�P��w�z���k���%/�^��A�k��d���hⰼ?W�=���<����E"���4��i���H#�':Eii�ܠm��7�*���01g� 3է���{ۺ���N���#+,?����1d�M��4�߯�wBN�DV�!�D~��-�UC������d�m+�OE�7 ��p�tL�ML�y.�Q�Mw�&��7�Pt�ĺ�3�e��v��Ƨx�]���{51UB�H�j�S7S/\��èQ�Y++�1z���x�>�mVR��s �TѼk&p;dO�hF?;z�_q���0E��v�H�i�ឝ�V�5����g9�g��������ZY���'��XL�������s9y�څ��ii����::�bD����xd3�J�gާc7?�� ���	�i�.���J�51�xZZ&1�Hn��a�:?��� ��Z;~bD�%�:5�N����^���Y�J0=65ҋ�/hnN�gs�L���#��eL|s2e�Z)���Y�跾�ž����p�Ǐc�~�~R����EE>vGH#z�tEV�9;;����!#Dh7�&"щ��j9\�ŊY�<S71��30�aP��s��Q�x-��(@���lP\(�� �m���rQ\W��VK����R���O�i2$�A��]��[�"O�S�mI�z|GY�[|�~�p9u�׈�7��?"�JvL�y�������Q.�}<Xm��]u�����{O��}�}" �mg�\�޲�ڲ��<�F�D$j��o}V�eWAxW+O�m����&��{<>j����l��tl�D�m�ږwL���ݥU���ӿ��Kd��y�?���]��2�*�ܜL"��N�͍�R.11��&����Sc��1~^�ͮ�jZ�\LӼ���"�!�|�RLK1mpO��	���#=�}����Ҵ"����Ғ)x�P��}��N6���v�9[�{�7�o���t��)�����z���w���I�x�T�Q+�/�/�^�:�Yl���ሒ؍:L�`���w����4/eIӌ)�/���QGdH�(~	2��M�=���pT]>T�'�
&=��<�Nk9X����G�1�ek®�����x	CY�N�;�K��G�����TM�
%g��*���Z���n�I@Sٍx�J����-�Ȑ9�Ɖ�k��l�.A�:~���,��3~c�"'����;���)18�Gï_��&a���w���<�"]-#%55<�r޷��/��� ���ԍ�ڬ��YM-fee�B������ٙS�;��ˉ�X���䏪NqF!ըT�r$ �� ��ٍ:�N���ΰ[uhݥ{�!�*M[�>�J�;����>C�[���{ȵ�޴o����>�٨Ϯ��j�[�|>*��z��gdq�L)�@�7S�o	P����߭^30G��kIER������,���Ѷ�V,��	���qMO�C����)��
w�fP���4㹏���JI��C��<H��|r��6^�e5	A���gw,<%�By3��qe�H��]C��\��W�f�U��&=g�t;Si�%�|��A]����8���h1^Q��s� ��ϖY���FO��++3,�C�����f�E$j�7�[/+�M*gMFf�L��ޯt��lG3�D��+�ǫx���)]���f��!%m^p��ƯK+�����¶y^X�����+�����9'��Tױ��kTii���+r�����ʙ�Y1z���J�,�������퍍�^�9��o=�Fd��<�|oo�F9
t��
���kʊ�4�\�@�l� ����3�ш]g	$3��erG�*�?��u�M�.�L?�k#A5	S5)�G�:n��T�b���
Y��J=Y�����5�	������nx"�G���T��i�dy�����hW�`{t�pl�գ�"EvuH�oT�/�g�rt}y .�3Qz�&9�77w']cF'��K*JX�m��3��T~�����!ÕT�j��F{� �Mb=<�b��ė��6�C��y�?.��x�<>>���_���x�J���e�E���� "���/����ļ�,U��V����S�]�X���4"��/_(��`��ه����)����+��瓎݅���*��Z���D�Ǯ��" JgW�[M1�����>��SN]GQQX�ߕ���WЎ�ͲM@m�HV��z,
��+��y��R�7����#>8��P�#��9fQ;>?�0l�\������t�+�)�\��h�I@ZM����o�{����_^vp)�?�My����S���!_RP����h}�^������ֲ��2�*-��Ɂm�& �'����7V	���y�����ƒ 4Ԑm���<C�q��)�W�A�M�>��m�_�|�����Pؠ�*�cm�K�	�w���A�r�us�x�8/�X�����b���߾_Ŏ�&=:;��WT����6n��w򶢫ag�c��XZV�N��S����Wf*��XR�3 ާϦxy3�j��`��Hש)������],WVV&:�	�:�Y��p�u���S��F�ǞH[�<'�s�K��m�|��bƎ��`$A��	p��%'�"Pۼ�4ʧI:Tq%$�f+̥5\��Z��r��V��B�{����*c����~�&�mi�v��b�`
	�g��xa�)�)Ϸ���q��M쁡{qW���������*Jì5����J>����g�Y$��Ic��Ų�ܟ��WϢ���]p}�gyb���4�3_Xv�&�5��뾵��}?Y�\/��|�"�w��f{��6浶F�dQ�Kt�RU�^�`�_�8U�I�BB�-GNir�>g�aώD��D�y�L&&�ca"�}����	a��
�5πpo�?�Գ�����9��g�:�gX���v@ۀY�be|aZZ�� �氏��J9cGmm�1�	)v<s�^m�t��ƯMg&?����K��/)�N�r�rn��SB�@�B�g��y�����l�+�s���0$=S)�dfg^���`����;}l0��4ة��u	��m�����zi�U��v��^J/�8��t!D�Y��tZ���{"4k'K,HuE�z��_�����+�{���R��h����U��}�ӣc�2p�Rn�4
�"Q.{������X#B4�w��f�a�ۇ�/N �7�N� ���eYO���$F8̋���2�WTT���U7�xu���}aa��k=d����-R8��A�f�>��W�'�n'J���hm��.G3��6K��:dd���'ǽV����L%�\�p����?6i�鍁粌�7Ɍ~&�S��r�����Y��[h:)g ��|'�G�n�j�j.k?<S[C*��~{��N���q�#+�&v�]�j[Wp�$tΖ�u�zhp�7ѵBnf����@lxI��� �7���D�RD!���^�kM����[T^����Vј�٘Ø�������	}�ħ_Y���lzrL����6�*� dee�?T����:�G��m��/�w�n.a,����v^��D�6��j��EM���7�a���.�$��Z���Aש9���6(�7��$Ɍ��ojTO�@���^��T�j�۰/6���W��f�!؃VSG�̉JA�~HtƤs�g��]�R�@�Q	���8�~���D��1&�x�[���!k��Z@�`T��n���^�crrQ����%���Հ*���3$�"� ���^.@\�w�3��n�'�<ڽv
h���Jo����&� �ؾ�~�o&��{�}����I����)&��x������Wb�By;�{�c*��(��=�ÜFݯ �b����E�E�c$C�O`H���iM�o�r�E��
�ԏ5��<.��Kl'�(T33�,C��N��uK��9;V��T�ls�k-�Ae��7'�u�k�m��W�2ԩ�WL#��\����q###�.�ﲽ���x9�&�~^nNhi���,������va����8�!C�3�����-"&m�L��Р�F�F��[��x�S{C��W��U�,e��5�O����E��B��J������zCI���45��u&X��o�@!'�Eix#��e�"'G�����b���珲q����=�a�����ay�$�f�	��s����̐b@����q�<c�S�3�(E��Gﴕ��]6�ׄ���~�{h�ߑV�P��)��Z���҇�v��|��j�܀or�[\~K�ڳ�����dUv���6�w@;Oԙd`rf��K�K�ea3刭���H�6ϩ�%��E$X8-.���P��i4Ql�a����٫�WX��ߓ���kG'��jg�����Y�I��ԒީaxOwL��������ث+k���( ��ﱆ�����sul[�LG��r��d9w�8Ey�ڲU�	h)�������59}�QR�B����v�#6�7���W/�d��V6��6�$NF�ާ����>�.NMY��;�׾� N\N���2\��O�t8f��3&��-Rj�<_Jtܯ�<�����H��[�1H� ��_E�//+;;;ǂ�FG5�Lzx��G�q"��w�=�~�z�PA���[u��զ�r�h�s���͂��:�@���jh~W�{g �)����\J����(vkŗ�O�~Cnx�pqFo*]3ϖ
�m�ȮS�X(�#C�1?�jL.{H�P����-9��FԊ [��CQ,7;���;�G�V���*�~��L��yI}z�e���	I���
�E�ʚ�����g7��Mbp�3��tâFm���#�y�x;zIi+���2`į�E��z�I���0@����-�
SX�BR�} �R��f�@])<��*����0���s�;�g�j̩��5��&��:��D$�~�.�O��i���� ��F��/�0�������+̓���&q�㿿�2֔���Y�8x-�|�����q�ޓ �AG^=�|I9M�2 ]��^������S����	؜ ��R�R��gj����~��uu����f��@��Fs�r5��BGmz̹�7?KK���@&"{{�7dQ%B�@�I����2׊���.Lt���!�7V�����_�{�g�s��1��j�&<:ŉւ����t_齸���b���]�y�[�w�m���zuJ�Zȩ3�Ķ��]Wx�h#X$�S{� �L�oz��AoU�K��tP%=���I<��,��	O
?��Ȕniiy�3g��0�:@��>�����Ne�]�����k[���9]��?��.���geۉ�����A��w�x�7kʉ?cћ���S�L��1 J���Z0�PMn
�O�kؿ/Ք�O��uY̔��UKn���|�r3r������a���icr{Pw�±s��$��鳅a���ٯB#W�[^\X��?����"�:�u����b�[�θ3����K�s��&����,te�@N:x�9~��Vsp��!��8๬�u��}�Y��l�I�H��dm���Q%2��>���&)���W��Q�����5�>Z-	���"Y9+a{݌��@lD}����F�:o}b�����
����7Do蹢j�vPD�NP���aWEU�L�H���o:��\�>f�R#�<��j����7l`1����w��w��6��Wb;=�;�K�t �Ɨ��ҁ��Y���?�"kK��z�.a��o�M\YYəZ�\ �RSVr�jI�T��V���C*�ڲ �iޢU P��:e.�\����Ǘ�m�q�?{S%vN�)F�6^�u�G�j�LOB�o�?ηo���0,�IډO9���ņP�� �-7��p\^�r$0�'椂�`�3�}�.k,���'��'?˪�KJ^&�8:��\����� bff^:��%���EJ�5�&!!Ҟk|U�f��ՠ��*�\����R��
�f���3�v��utd��i�8�h2�7�Z�7�]��R&짛�A��5��w���>��������z�5f+'��r(�x2�8�r^.�L�"G�

�UR��a�f���x;t�~�)
����-�&�\$����r����B���_?�A����{'���hd�!,��X�+�Җ6��2�rw�V���5�QxU/�ŕ��IUu�݌��1u)Q���[�l)�D�B����C�����ͯQ�Ρz%*���B;͌@mM��l���vJ�K���s@_2��)}}}��M�{���G��vS�!b�&ݩ��Y3e�p����B�IK-B$sxg�t~2v4�.f
8-��[����z{4�����2�DF��/OY2ʉ���b�ֶV�ϟ�������j���&�D�㵘��h��C�4�����q�Q�F�gF���V�Յ )�z.PN�H=�+-�HX��y�ru$A+/t�w]�zyk�����A�Xm:�7� �Ӏ�"�@F�ל�~����U���ۿ@��ࡂS����'4H��M��$��spm�z�w�y`�'1�`�]�q1�n�ĸ"5�� ��֝��z:@����d�jh�u:2ԭ>_w��ڌ󹸘kيse�9>׈iKS�m0@VJ�1�'3=��w���$"��"{,����F���t���^&Y��T+�+g�k���#5c�e���Db��?��é~L�W����?fSjJ�i�JH��K�Rf%0#�{�n;*���}�~���N�2�Q_�S�®L�Q�qG�2�>�O�غ`U\�ۉ����<ި{��<�TWS�����%��P��5Qr�Zc�ǫAيE�_�"CD�|���|�l��9%k9tґ�?����
tȼ�����6��k3�ҭy���,G��� ��9����(׫.Fry]Ͼ���a�kJ�����PPN��9�Wx茕��pJ9 y�{f]��i��8�1��`���ۿ�*-G�Pq�(L���o���������.Cy'�E<[�/��O[%�	"����s
��I<�)� s��(z�'�Iu���8Q�����J�aI'�bĉ�u�(}� ��.���p0����BƝia��� <\�r�dc���#.������yAM�Y���X>FW��$~2iţ���2߷Ha�r_�9V"Q���;b�����E&_w���]T��敦�ǵ�hE��Dk��wHc��4�u0�Gɴ���� x;l��B�نu%��͙
UI���n�֑��V�JuF��C>�7��G�-�+�|�D��n..�	?�P�4����s����3��Ս(�º K�N�,����g���c��7�$fɯ���r��v��펜�{�8K454�d��b��ɰ���ws�>�@XD�s����2V��$S��=|�舞2JCW7v&u	ԩ������烵Yd=T.J�jC����L����X������m��#�����Xt�n�H���t�Z�d�G��@ l��ss��>-sq.dG�'�*�z���+�"��s����,�i��Y8��� �%l[4��߬ۦACKK�'�G;M��U���6\��G:�=q���/!2]����W��"��' ��ʊ�Hc���}'+u�bY�����n)}�m����)$_5v�V�G���'6w�b�9�U�B5�&��̞pd��5����'"s74_e����;v"�%}p��r6*�]�ł��aot���	�����"ߘ�Ŋ$xE�d}dc��B��R����R�+��{��Գ����.!��SK�K�g5��EE-74g�`-*����9Lӓ3o&Vւ��+W�f�m̓�;'�V�L}QUˣŋt�b���{c�2��|&�1��V[~kk�����:H�yl�L]�0��X�k0�I�k��V<��?��������{�#�k����m��H�;�׹<���p�<���JNM��ؓ��֭3>���̜W���9x��qAP���Ej�
(�����	���C�*xVnog]�Rm�g��POoYq��o`bo�I爑s���	�C{3���nN�(�����_Za�5X9a�3�8����`Oz]^L��ͻse����3tZ��HN-叝Ί>�<���1`��;�����l�D�@�]�������xdٟ�߿���p�&��k�ׁ�ϯso��h��H���@a֢�s���uo�z#���?T������{e���UK���.��r/ �Z&�::)��),���gT���,^���у��U���8_�n�����_[�W�Q���^�����h��?�}�H,=�9A���hVW��T�#�쀁I18{e%rw��/�w�唔!r�ֻ�S�Z}������Y]�H�K��Gʑ�#	�b����@:��	9-DO�B�ɛ#����w/������1�ꁞ�܀��EާgiQT�x�#���������R��~�C��f!�c;�zDa��}�z�Rɛ�?Y\Rd��������](1n�\����(z@�����&`���ޅ��a.s�a�"�J|<�:�p�Ov���E��ݩ����qV��@ZtV��� 9	ϯ�8������s''&2�[�g`�F7+��`v�����F���he�>��|/!���U���������'kC>s����\Bz� ��ĨfH͘��Ѫc��������ӌ�Ç��4��͏�]]o�4�,K}�O�枞j����.A���-���x��:��=Is^��OI7�r�i��EEV` h@TM):P����j�E�kk�m�''4��>�)���Qp_��n�T��M���?��o�pEGwF����)�8���	.
K:��M7�ӈ;�N���"7�qP�@AE5��D��g[�U7%sȊ#��B1*Xm���}���0:�|�gdb�@���[ssI-O�ֶ�)��y��ăo&d������R'�����8;]E����+t�����?oL)![K�l���Ӽ~c��^�_Ơ�9��DS۪�+e�*Q*Ƶ�|�W�j�\�
���Uk?��a�	f��b���L ��?7X��k�xa���r� ~�K������;/W��x��;���QRo�>�P����"�"��yS��1̏g $chQ�¡�<�U��<5�Q�	�дB�8|��̀�Y�{򂷶��eܩ:�;�H�ߌޟ��lx�]nRnt�����"�*ݴ����b���Q��4�R���+o��K���h��i@g��L,��m}��L��^LoK��ag�م���?k��yD�;eS���+��0n�O:^Y��sK($%%u��"ۺ�q (ᠣ )���uٛ���˒ϊ��俣�o٦q`kL�
[�R�j�*��^jJ��l�pL'��m��"�e#�*hr:ۤz��,-�ﭛ�B�DD�^u��g��js*�	�O�xO����6r&J�i�K��:�QC��F��܅Z~����f-1����|&u�B����f�]J�۫L�tuw���G�U�E�|}EJZR$钮�E���[BD�vY�p鐒V:���k�|/����{���ęO�9sY�[\/�����F�~��!Y���K3��q��ٶn}ݔ������埡�w���\� &LL��g����~ ��{�^�,k��Ť�L���n��/���5.��fû�11��p�C�R�o�R�Y�ڤ�;���y�TxX���n�y%1�\�k�Z��(,w�f\��y�'�	��Ϲ�4߲�K�=j���D���f��� ��������~ْ��=��%������@�����M�]�h�U��AN:5-�X������{
ŉ�=�]艊��jl�S�7C���z�Я�$��F�`I/O{/?@ @����JL��!U:�H�s�f������Ԁ~?ڙo�yg��P]�VUW������d�8��FXܜXxl�666���?��w�!����b�p�{i4�T����O'��)��-Z��ݚ�����a�r�("�apv`~vV�?�ҽ�^2FD�����m�F�XI�~k��S[�}n#���N�]���ȒD@H��ų��zA+&�#zE��6%/���i��i�ltr���y���N��?�l$���#'�kg�j��G�<�la6��L�|y������uL��4sn?�q�c��M5]��[�sfh��_��-L:h��|�,J��z�m$�ћam�4'�Nj�=���ݜC�7��=Fg<B���(�|{�N�.ݘ�R�K�K1�׿�|�EŐY��j���Ǐ�l>��(((RRSu,,L��Ib��-��)$��Ӆ`�!�R@i�����e)-T��KLE��״����u�^'H� �Ю�:'Ԛ�P�TY�4�[���
�c�&�q���6�SRӴtu#�-�W�~���9d��_�]n[2{5
�>>&����ְ\����K������\vԦL��ˎ�R��������c��{XN!k(��8P�%�C# @V��� �Ɋ�J�Bk�h��}���ب·n���~�~`��mr�m��d���ϓ���,�aAG��(*�e��eey��1�%�>��-6��ϕ��^��'��B�	�����܃A�����el���r��W+u��>�����z��6��n�%���ә��"G� 4h��q#�"�%h�S����խ�f�J)��r��H�0�e�j
늒��Tq�O�Q�~���*���+�AO�F�՜�{��f��0���sX�5*�UIs�}�t���gkjm�����aR����{���Q���ƕ(ɬc��n\�����Z}n�P��8�*�1���1ԕ�"U�?.AXh���5�6���n�~sO��M�%�[�ݤ��L���bݻ^ޤ��p^��m{f_�$�����X٤��/�AB����K7r#%�}r���R�Ҙ�:��d��O`�5W>�F�$����j���uy���n�BO�������RV��/�bm�����/E�*rf
wc���\�gƠ]��K���0Z��-��"zUZ0eeH0�E�WV�Mb�~9�U~Ƃ�L�!M��b�N��Խ�F���#H�I3_ɂ �m� �&���hU�ޡ �r��.�U8Q�p/� .J&Z<�B�Vx��R;Ky�D�zEӞx��]DCf8���nAUUL��4|�e�vlz��jܮԨ�����o�)���	��b��s�BBA֬�0���rY^ϊ�:j����r�:TE+��R���.s�Ն�OQx��J���� �,���-��lg���͟Z��*�w_�|�ӈG8dq������s�&�����&	#Z����,�=��-�������8*�zҩ>�����@.?��_�]akŎ�U�����N�$��Ą����$?�k����4���ΜT���c`?JMU��A�V�-Ed���#���l<��Ctx����L���������tC:�Z�n��7?��E�w6�?)�(e��I��Ǝ�����W�T����L�EgL�xxn.|ܱ{_�cJ�X�N��U�U�ꘈ�K���ꎪo�[=аiJʟ�SE��?��1"����P���~���9R�HIKc��q&�O�;VL474�4l��K0�pz��`�<���ťi���`���)a�hhht�+J�u��#`�gFFfA��14����hKkP?��4ODPHS[;�i��1Ԅ��t)IO�����(	0�H7Y`7#��0�k����L���P���C��-���k%t��=���dN�'TM>�NN��MR���wP�[�$�~��GHB������Z��;��[�Xm�u�~� �`\�⃟��O	{��ⅻZ�>�b��^�P}�nV��� �2 ��At>�ݬ/؟����������˧�6�J2쾾����w�r�	�8s�����?���k�>�a�}�\����/)nyJ�Y|�������H�*8���/�p�^�	:�2}NP����{)"��%J*��C�?y^Y��V�>�@�������zBm2��<h=�`p���7�+���K��`�eD�yaz���-�k���C�۟�/T饂>�UW٣b�o�A�c���*�h`Ľ_?"�ע�i�<��v����K�ؙmK��+Ƅ"T�~K�.�w5\�>�ANE1 B	����?�[�������fgg�l��x�U�σ̧o|�L�V<����\�G�K�/�����楯����t���f�]��ؚo�SOHV�Q�,A������̖�il��]:�rN�R����IQ��GF��Q��e��w�aS���-<��9 6˧bV��R�]��,:O��\v���sD۠x_8;
N}�Z�y2x� $+(`��O��Kx��X#����22<�Sl��9�R�1��'��O�iQ,/�����B���	I���A���W�boW����xKh���Wg�x�G鶕̺�p!���M����|T�tƪ2�2"O��f�3�RWI�ZMc'/;�;���ߨÆ��m_]kw�/�/q:���KlCcSW�{��#5S���<�nǬ���I������Z��B�Ή�Q�	�$��#�ZZ|�8�x���Q�V&M_c��7�&�݂�|��F��f���o9�j=�t��,�������ԝER�):�8��v����#ܔ��+4���j��ߛ�>s�ԅ3�/ٻp:�F�vk�#��������{�/b�1����?�F,�CT�9��9.zLe5R��Vf��vd�sp��1)s�%���s������?ↄ������f�=�uf����%Fc2jĎ!�9\&��W�����-�ʩ�Pt��ibL���@��.^ý*x$��13����N͍&k�b�hΫ�g��y��)(8����!~I5�3���ts���s��_5Վ��B�Q����{'*�� �V��k�*��� ���``n��L����������x����1�<�j΍�u��/�-��+�>U��|�������]��/(��l}0f�����VJJZ	ǔ�Y��7M]mU,F����ݎ�0��:���������
��d8�;_`]]����5�bS#�O��P�lSIà���<]-t�@׵\�1�*՜�N��*_A��qQ�7���ht>�=��PffȒĊmHF��rTܱ���`s7������>yb�����%&�VVQ��`X����5��ƭ�����zu�Q'���#-��QQ�;-�?<�疩N�f��o!��u'�����!�7��J��y�k���t��9 �x�E�w�5=7���#�_�fQ"Tl�Ռ��Q��Y��H��_M���1$���!���x26n��W�䛈�ja>I�,�T��A<��b7�#���ˊqbE�6M+���z��l�#㺎��K��qG>���<�+�~�[0�?�q� _��!��{����ʬq�į�#Q�]~��
	����E���x���3�,=�C�P�����r����}wʦ����v3���VH��R6�N�&a5�à��B�I��W<@�,�҇�Y!�MG���)��W�|������ ��j�ڤ��MA=G���(���fiI	y"L)�gy�qE˺1 �8�Yi��R�� K�z�5����0��)ݏ�J�M==�_����Gຎ�����(V����m-!Aok���A��do�����\r���R���������6<9=.�-�l}VgKx!?��ȋ�q���Q�z� L�y�q�kC�[NC��<�ddN�G~���C��N�\���]m��5��F����W�@�C�aS��̵�=<-Q�AvB��Uǳ���zN�ǜ�pG�x����{Z>��gzZ�����q�Yr�뷅�. �.
NT�z�����_Τy�GP�nc�qZ���Rv/R/h*u~���!�qq|�k$y���*�Փ@��7C����oRd�7��I���|�I���5! ��Q�t�q����>1��
:�����!�G���d��#Qh>~��0/�'t���zzG�U�<p4iҥ-��V��vW�0�[�fX�œw�g�Q�2��㢽'��*��P��,,��gt%�<�p{??�K���4}5�Уb�(���;Ya_@��X[�A�AU\vC�4�'�_��q�W�QC/�w����䌔�����%��UT� �����T�"��nt՗���WU������|�͸��P�GϷJ}�]������ �,�R�D�����t<��$c�6�"�uҼ�{��S�'j���.z%�	����zY�̋����o>��	��"n`W�u��|O�sJ_:j;�3�>����s�D ����;�^\(�dG�a��[[,�i�GN���[�1�,�?c�M���>IO���Z�
ND/^�ީNb�K")�U��{�o�s���I�t�R�M�A5]�*뷞&K�D1$e���6�j2ft5<�E�~8�$	E��M2[U����Y/��@L�ʊ/:d#�?*i�v������V<l)��2233{����*����͙����
�O�STQ�WQQ�A6EgL���/�6�����Z55a�?��c��P�/��<�g���+�]725��d�Tr���NbccC����@��<qǴ�[�������RZ{��;�ݶ� �D@0$��iu�!���LgN���D��r�y}W��Q�w�BM�8��m�AccSQI���
~<�o~�9��'$���bdjl�ngm�?v�mk�8}�:uhMJ9���O=��(�(Yޖ�e6�dBmn��wр��ґ��$I����9���A�ڂ6I$o��֙赧���5��
n��u�بY��̄[���S(H����b?�Kr\�L*V[ea)��YW���>Kې����m�����\w�Y7������?*�h�,���W��jK�&l����5~�����y~$�wj� �WQ�`l[��y�;�D`�m,��������1�%�o��<�{?Yk����<�`v^���ש34%��x���Te!�ମ�vX��%H�y5u���}�G�)���3��%��iˆ��N�}/�&^!�U[���o��/�0L;�~�m��/A�D�L�!��C.u����s��&1orq=>TW��3P�/"�)��g������`� �H
��x^�}Z�ˮ1�%4uru����i`�~~~h�#��skgyN�����0�jQ7 �
���(�g��2�������i@�#����Len��ç���t#�,��~�-�L�-V?�;
kk��-��>�O-5ӥ��ί�$z�XI����h�nr�c}�u�p�C칩4��JRr���JS��ߧk!�ˑR�n���vY���î�/��L�i�rZa[[�2 Ʈ��l-�X�"����8#�I	�6���� �ed���I�s����^*��g�\;.�rlM4���'ޝ�!h��<Dӯ�>b{�)�Er�H/̙�\|db�v^�Kf�̈́\�`���Y쐶�sk+j��7j&ZS�ÿA�2��<b�(�={f��{w�q��O��g��Ml���-�����6��qe3�,g��V��#DIG�CS��ר?X��x[�I��A}������E�4�s��ݜ�y�����]y�򊍤�f��BB������~6�r{65ג1R�I�f� $�'���g��q7*>������c�D�{�ƥ�8̓��R���S�K	��3%H�kC�W��7��
~qkn���;]�EcA!��������AH�i�5f|� ��rl��t�!���rJ���aàb&����i�4����Q�?<]<�G�haf�*�*�lM��F�����A�=�8x� B� �8{�ͣ!�����+�J!Ғ�&߲!��ciiiS5��*�̃������	���^����.Hu#�^�.-w� <&�3%u�!ӿ��to1�U���!���ё�����;�W�ak$)�/V]���	o+p��-Uw�&R��j 2s=5�z3�J;�cM���O٩TZ���y�2U�Jm�6 멲�3�̦aj�������-�2:^X��7�	d_	����7���QMf��%���H$r˂D+B���h]�S��qzb��$���J�m*��7�������O���6�c�7���U�R���2�~��=�z�z��侷#�&�>27�����C���2/ܞf�	�ˀ������.��-r~��WN��z��++t-�� �"r�=
�����m�d���L56y�C,uli��ý��b
������������C�Od!��`�������� 6�+W8Ze}�#��FC��Ad����܌�����YYku�[}�!Y�Ȧ�?���$��)^@�O��2�bT�K����������P�>��Y��ϻD�~�m���]���
qk�7�h�ZJ��{� I\B�9���,��r�]�v}��~�㶭$�����ʌS�ޜ[a�,�ł[�K&/��\���ys.���<V޽���qK=�-$FQ��/�4k=�c��b��Cc�1��I�;WE�~!��i���8�Мdۡ�T �,��"���]C���;�<-�G/ȹ��%����h��kvȌY�ɵ'K�/"���S!���c�Ji��{�ii��v��H��_�R��ý%7�>4"P�Hp�����;�j��k�)��&�:��*�����`�dCl(M::cGD��^ʚ���u�ˢ�����H��k9�/���g�eeg��Af\-��G��=_�*����ed.�1	�`q�{���X����	,���y�d�:O\(����m,�4���M	��Þ�N��N�D�M���h2�lnh袸�pB��1�+�Y]
g�[߹0��﮶��s#�Bx���x7q�AgW���p��7��+�0/x����v��w�g�Wqy�d�*��.�!-\M�ޞ�X��g���{�X�?��d���f�9���ݿ?�IN~,��uX����3拍c1'��]�OkOI���ެ�o�V?����bs�'Ϳ�v��p�2ݾ��k�M�?���N���B��Χk��#\y��L�������]w��6&�5J6R~��uVP�v���J��LN}�Qfd�(.�B��˫Q�mR99:<���I:2�x=��C@H�r����j �\�b<j<"�7���2�yb��d�HI�����		^,�
vj�8#�&<��r«��6-�����D\��6?/�,emc�>������Ϭ���3��t��;n�}|Fl�ō�pA�4jǮ�8��Gxq�f�[_�-\�.:ϩxl����.5�s"�P46����L�$�r���++k�!9E1ǔ̵��"4�-��̬{�P�� n�}^eeB��c����P4�b�K�־A�f�I\����%QtFF�Wo����iʻ�"�6WB��F���X��N�V�B����6��]�Sg �oW#���<��y���:š�H+�vb��� �9�<�y�>_���r���*�^1���� ��tהq�J`i�ѐ�gm8S���
����?h�y����Y�LR2R��ꑑ���us: +fgUj�X�����2?|>�7��|KJJ��U�I�Q�!�����g"�os�Uu������������z�64,
;���16���gd�m�ϙ�Ըv�T�L����;�'*�����3^�{A���&�+�hؠ�*�_�eO�غ��u��v5r��[�!��O*���ZY���+_\������>LK�<�ቦ�:
C��򈉉уnA��`)	������vU���ݽ����5�w8X������U�N���s��������u@�rrrR/]7�`kSU+�e'�����zN4��LN
>
��`Jж�*��Xr�Z���P���zh��67s�'-���k��t#M�����	G���Sr9�,P�_bC��BS��/ي��z��X��N��	��Iҗ
������֖L�Z�t�Z����Y@!��t(�+��|��F�r���p�A��tt���i'v˲��r>Z/i0�#��j�G�?G�G��xW��=�0}|T�A�t�Vj_��*	�+����o�����˄�K���34.�5nNX=���";$>����~{�\��W�8�
�["=�rʗ&��v�B�㦁�p<�:u�����G#4Ϟܫ]2�=33N�K��wh�>;��+��iT^�J�#B9q�Ua�Q�X{��<z��8�������DS�$d��jQ�-g�e�S��6cK��O�y5Ȇ���)���޻�^�����I˘�@0����X�3���l��L��9f�6O��A����Cٗ�:~�����z��.���4��F%(ڗXґ��������d�W7@�HE[\/�2C-�';�������S�[�˪FTоԟ�)g�V����s�I��x�ɔ�=헊����ch%J)
]}+}����@RN�MW�I����6��N������_H����P�����v�}m�ƛ�eV��b�x��4V<
���[0�����%E�;�Bąa�8&]ٺ.Vx�ڟ�4�_I��[c�-~��7�Ζ8���gv���94Ee �oZuEm~TSS�Ujy��'����A��\�5����V�x��^���½ռ��V_��C��H4��| 5I�\��
�>�~��N���c4(.�ʗf����O��v��P���x98�,����p#2Y�6��-�̭gӨ8\��Ȕ��F��:\H��a�$#�����j���K\��GEAQ�V�w	Z8����X����_��j ���Z��ѾЛ��aPr6��g�j�R�0��Y/���I[�t0&^G.�c���覧���C6��:�ó�f��N���h�{���N�Q{	tr��	.��\)��NC#��tu�G�E����P'��>��Cge��d"����X��]�H>HP�0��d�f�B�^q��]�����ﶴ�O�*��k����^*a�de��x��DS6���쿇1��yuu���Y@��+2�HvD��������c?2{�ۏ�Dm�'C�mѬ�kX Gt%�4y�`\��{�~��B*}Ӵ���f\��L0���ټϊv��ӄ�����7.'d�-�	�A�d���#eCڲc<��O%���}^>[Z�n�;^j��˳�����cb�5F ���{�81���TPP���A��D��H���?��u&N�v68�	i|�3%ac���evw}�=��e7���GMDjjj�#<vc�a/����h���l����� ���Y���aGGx�U~`���H�(W��'���(7wwm<��͍M�SDxQ�]�ƅ�²2�ቐ�N4�p5���L������Ӫꩭ�mLB��$�bW �R�/�g0�$�����W켼���j�>� �r��fF>����~�h&��^���E���lx���9���_�\vy��^�h�ܘ?����P�r�#�/-t��1�}.%�żc�^�^b8�^�E����$�ddBm��({�G��+FR��?��,*)��+�џ�"!�p�Y%��E�&+_�-uF������g[={E2Hen��>�n���R�+Y㈈&f6:��o�-��?���d�s�d:L���Um?4��u�]����)�D8U�<��V��A��w$-�'�������x�&O���־ ��;�%{�5|L��9$&u�̼���%j���e�<��~�MHu��]"�x��zӊ��%����!ڵ2���PQhT�_ٶ�J�{���h�J
��W����^�
��0U���d��c' cE^4�W��9��|���~_E����$�g;;\�n�%%Kb�EE�P%�&Z��bm��l����ߟ<sp;`�Q���H�S�7�=�T�~{�k2�z2`v=a��V�ccwq�ؑ�)J�����6��� ����Ed�=�ٖ:ivft	�WGbo��e���<YbW��!��[A96v�p�p��F-Z�+���/�ii�@�n/.V�*˷�X�������x�Nb߆�����Z�n?|�rr��0���;��<aH���8r)PF)��LT�,��D�n��z�}�ȗ�Te�RL*��gf�-W}S}Ȫ�>���P]�g�Uk�+�;�-����~�4��|GGq�8G#��͐���m��a�Z[�����f+.�AZ��"EВ�R�M8�I���]<��J^􌡏ʱ��2A�A�Ӽ	�mF9��AUa��z\������3���7Yr��M�_#� ꯀ Bj������Y<i��W���QVQ�{J �T���g��}z"�+WLnY�ǳƳSp�t�=^���i�\`�+��r˚UO^=������\9�Y���^�z-���ak�O#x�-X�,tY
ZV1>����u�2pC��xx�I/��O�x6���P(�^��Ê�=�q���S��e!�o�Z�@�*��m-_-��`e��{�L��r�}��í���T��zQYY���J�u$�Yh����T0N]�Ii�$����WJ���vU�M���j-��!�Ӡ�l[��P#DN��㝍�9���ٍVԮ�1pk&bupp�/*����xz�3�4f���xݟkp2ӸL
~�=�����������s���$��}H0?��z�x�7�%$�1�]�
"h��Z
����77D���<��S���c;�aAA��R��cRq_&T�q�R�犃�^������>�%�_P�Zz;yV��_J��-n����Wf˼i?wB�ػ\_��)�d������%�}����>$�}����|�!�7�7����E�'tR���mѓ0��O��JG_p0,n�Lpj��eT�/����^�omm�f[�L�5*U��hh~��OϏOGu.i:ǩ�A5���7m�W��("'����21Hg�����3������@���������ƿ�<����n]}�$�3m��Q�p��{[�4�,zT���l���[�����`pM��_���*`|ʸ���wӀS���;�b�������Gxř���|A�ڳ퓀ړ�������#s�7t7��v��c����J&��l����|r9��{w�,�+G�ǋK,�[����Y�{J���ģmj�Y������M vw�(�^<IKK+��=<:*/Jkg��=�سi��܁�fk��� ��R3�xpS����6������-�uu	�l#c�T�)q���+�eG�F�l섍>��d������WVֹ�$��Z?d4�����.������ZƔdm%���|��|�FD��x�q��Y��T�k�Bm�ٮ�l'��fH��!+:ׅ:5ӾKύdIl/����0�nc����� ����_v��`�/|�~��.l��9QMJ�u�b�t����ȿ������n��8�y����^U�w�������A2�<�;��/�����7�t��D�i��ɝ��k7�o檶O������ ����<���[����m.��d�	�,]�^�~ilWVQ�y�t:e�|sjS둥ޓ�mx�j�cG�x��ct��,R�� ��w������SE������v)��kQڴ�v�����KF���5Ӻ\M�}"'?,$*�#*i�;00z���~��&۱���g���=�Q�Sږ�.~A@)c��� #![)�����.��Xyq�չ�O��0����j�.��O��m�*�+0.i�� �KH4�C�$U�ԙg�pЦ1|m͖ [c�{:	O��UH���G���=a�h��Ӿ��r�6�6llr�q������0s6��1rJ��H��.�C�O��<�tq�<k���6��4Y�f�Z���ֵ�qx�=\��>��)
�>1:}���VW���7�@�`V��������>�-8��]GP><7�!���� �s{v~-z���D��b�C� g6��ƴ�Z��|�E6������;�g}Û�*�`�,(y�_����<>�o����ޜL
pL�KH���O��;�4����/^�ȫv������������h�D|��/a�_���������p"J룦q�ov�/�I�#�$O�R��F���YKle�J275�����3��!��� �f2�xw���tꬵQX�(TJb�R����xO���]6��$���=����(`���\�Y�I�q뼔Z�J��J\\���aE��?���l��ҷ]d���S����hm�����.���G���V	)j����z��:j?�c��c��h��h�	�=v˶s�`��%*~|�Sb����_B���}Q��P�����<K::@+8��! �c�y����n{K��h^�W�ڐ��=��EP�ڂ)�K��CI���7�Ŀ��x��Ia"�\�s��C3J�F���%	�?�z�7Ѡ>Y�w�-�����v�	�F
ț���$Cmސ�a��������1�����Wu�t~ͦ�e�}�*Ԛ �*#�z�Ȅ����u����E��Fj4�Y� ��0�V��ǣ,��<�WϞ�mq�ed�-�G��e����<����YZ̍�����4u�d^>]�Yhfz�jg�&f��pT��hÅsn�캼fz�z{�.04N�����eb�9(j�S�{� ��P"�+H�v{�_�[���-�����~id-/����˝����z,�������?�VY��-e�����eE�?���o�,Z/(��W�ct���Ao�jC23��cF�{�{����,���i�4ѕ?cj����g�8�\^р����yr|L��q����gX�DO����P���c�k�[��9E��(88�:��w麪G4T�ى��a2���`�ҷW�gg������(��k���KVs ���DKK�y�y�AǢ�v1a��"������M7>z���pF��~��p®��X���|^��C�����Jo�T<h�^đք�0d�<ʾ;�>�H���y����� �eu�'{��	���兯Y��Q�s9O{�|� ��}���Xc.�9��;�8�N��������΋�\�Q�&ճ.R���6��7O͏�K'��
%����nHڳ��5O�>�p�50Pq�A���p��-w�+�#��/�r�5ٺ��q�a�D�)<|�Ë��(�n�>�_�0�.�����6M�@���s$��`=�D�K���餸�?��+�]]Y�H��
(������4?��Br�C�Xڎ��3��Ubz���R�]N=��G�+	�����{�WU�ۇ~�:����cW������:���#�0���}��_�Z��{b%SL� �����!7�I�C|��x�m�w�oQ�؈$*Q���za�6�m�y�C�`V��kff�����-���D��\l��¾T0��F�l�e�`�uϗ.�(/��\�M��������dVu���C�E� zVZ<�A�$��[@@���Y)���{�[�zE^ҵv*�~a��8��}�ma�\sR�ѰBL̬?j�A�;;�#''��B��!���Md}�g�:�/�����|��Ea*ey4��.?~������IV�'#��܄�,w��y�˭�cTԓ7�����
~Z����%=n� ��`���\�YX��-�Y��In����{N��v>��~b�����i�A��K��v���p�
ưF�z������1�w���<�q����# T:��r���/V;��=s��a��!{��X��/;Κ_I���>��-޽:���\�V�kE��2M-�*�s>r"�Z���ЄN\�{ݲ=�#(~8��)#��{�6��v�-N)������BI���P�����)Ő�����~-��w+NPI_u����/B$�W$pr��_ZR�8+�[ZkaG�xQ��|��*�A��U<��*
���q�Z�J7���3�L�h��E��g�̸���# y|����g�s|�P8w�w

�Yf�%����n�	d}I��.���6�^|�[�8�s (7z���j�0$K�����o�ɬb���y��s��`���m�Q1.��_k��w	#��S[���a�r�	G^ ��#��������租�<����l�{n|R�sf���ࠤ�;~����DVIX���2ș��u:�E���H�)5\Ą�n�̿���0}$����O�nL�W�T|��$�qQ�L_o���m[�vp#⦹w�Y���?�R-nS]\�P��e�W���<�	���2H"hȔ����2�픘�?�N7�Uذӑ��Bl�'ȫP �?PPP����)���uZ�VFwn���E�$v�t'��%����G��q�;�����I�fAיY��.�%{u��]d�6�W���(`_?�!�4�i�E��ÉUݱ���k���0�-���^�h��CC���:dQ���l��ݨ�'DQ��{�'��w��qKgW��\6�o_\�g;U6�����eW�cA%��M^�a�3^Ҷ�P�b�"U�yTA�Zf����k�>��2�U�%��# &$�#L�L��0�J���9h��&TCݘz�5"�n;nt� IN��r����jjKhG'.F%�d?�����΁L�������ٞ�q�p�@�Q?���!ژ�����\+,��Q�iy6z@��Ňz������=���Yh�.�p�Q �l��t�K�ΠƐ���|���N�j8[08��PUe[4�w:}pw�JCsjk�s5������c����7s����';�W�5���3ߛ.J7K�i��v��_�w�� ,���F�_Jg��Al�97�=���x	����tNd�q����OA�/�ڟ��z���ܾ;�>���TR/�[��Ҥ�i|�xg8����bH`���t��99ފ;G]����ȩ���׌Jn��c���� TCCC����}������-r����&� Ķ�C���y���Vf�g<a�Zxa� �s4q�xG��Y��m����*4>c�=�r[o� }mb ��Owptͭ�K?���c~�	��_N/�e/Q#�_���R<Y��ڱM��h0����l�kg��L5~k_X���6	���_�_\��_f��{�����(��d�L�O�j�M��hS�Vây9;3��
���c<l+	'Lq��o��li	���t�h��^�Lx�bj��y旒>m�x]wGEV��wz���J^-��?Q�Y_h*�`m.�==�pƴG��Sڨ�����ĳ0%�{j�lϬ�|v�����H9Y����9ߝ�AI�(wpM����p��	�V%����k�����G{[�M���Y�J�YL+t����m�/?4a��{��<Ȧ4TX?r��skV��P��R�.����Ra'��o�V��N4q6$ك�,���b~Q����o�J-���`��~�w���F�����Z�?�F�BoG��m�q��.��QB�%��PӾx�"]�>nIذã�\�j��}�L����r626���+��d�����)��A�V/��̈c������I�!��g44��h������QA��0މp/x�i�F��X#<�V�����wa�6>&F����*��Z����C��%켕��&K�O� raG4_7�SOI%X8��>I�e�U*᫞c�ᕥ�c�К�z5�崲�B@dn��LOcm)l��f��h�S85���s��}�;0"�y�G�����U�F �$��"u�'��v�6�kD upQ�����k�/������(�G�Uݜ�n�-�8ĭlm5x]T[5�C�垛l2���0i�̄#���!B'��$VI�HE�Kp7\FI���
K�,��r䦗��3vnn== �+Qb.�Q�'�B^	�Jb�{'���0Nn���:��dWa���#i[�Ф,X��%��X�xh�����q?����u�O����6����co�QT�}�������ȬZ�<�g}K�Z�%4�����ߓò���������6���Q['�w�cҲ37ץ���dՆ1��n�m#!�ːS�X��#�N]η�]r�w=�`��N�`!ބ�sH���܀�P�:��Q������ҍ�}FƧ�obEa���d�Vpc
<�i9''N���X���Ό�pL��4(�v��qI�� �߈�K�p��j޶k~nnn~,�¾�T>��D�\	��>8Տ덙cm�A�l�a���u�[����BßӤ�H���U��ؽ�og��rX�Gc��6�P�
֖�Ҹhzm��,Q��N-�z�����K(髆����?*�>��RSO��$$&^A_.]�#�ļ���$V���Z��bW�i���t�qQ=_�i����AZ�A������AJ		�X�A��kA����y�ܻ7�Μ��9����U��bZ�& ϟ�w�%�ٛ����ω1��DIww��W��'G��hԉݷ@`�ߟ.�����	�ϫ�lϲ^��������\�0����=����Ű�����VV1i�Jo���7ǖ<g��Ũ���|�#.��+^�VX���	j�߷C���111	Xls.{B��n��|�X��6���k�o�p�F�6bˉ���$�ET.g��.��v����\�ꏆN����#.+2:�	~��}����o/ѿVm���ӑ���!��\��]`�'S|YI��88on�n�k���8^++��>��¸��k��crs�HX]Q���qi�N�wo�7���+���
���ڲtن���Ea �N��.~>��%dU}4-SRRx��m�}r�$�n��U�����0`�^q��o�B�;:D�s��O
B��zws����H)ڕ|�X &?�{�����*�9�Tk�5�U�L��046�O���r{x'��Y,�**�>SXca+�<��vi_�f���p1�����]\�	���=z���-M{�~�k�������Pi�'WW��G����x��c�zT�o�Y ��m�	f���GGjw��Ҳ��HS�D�����|Q˫�����X*�_��*JZK��Ce�f���N���?��r���W����$��V�88S++U����P����=m|���c���P�=Zi*�0%�Q}X9��w8~ޓ,�ҋ�虫Q��ӳ/�bdT]�`�J�)���zMu��ờ���9��dĂ�?|D��8	��q�H���b	$��Q�7yQ+��|8�@z��X��P�|�uQ[ŷ����F�?�ԟF�gB@��eT�C�
��b0��d�����3��ڳ�S�-�\���wW���K�s��������E�CN}�;��#Pzl��ߎ΁�*��9	$a,��Bv�u����õ�����  ��[�o'�[fNδ�C3Z�ϋ��24�{�腀U���0��G��,�1))�]S2�Ȋx�'����u��?��c�S
efe��T%������"�`�x�������Z�cUw嗳�RV�c���KN��4G�X���S{nɟՎ���_�j��8_A5O[Ȋ��R�N���9�DUu�W;���)��(�-�9��ߢa���Zԓ֤��yT��#A�ΗD)Z�3\l��u�Y����d�C�ɘ����A��h�HKG�;x�Yr}��TK�V?�r����������3����Z��rI��˫��� κ��ٔZ#��!�/��v���8���uΊ�;88\^_M�v�yTl����e���+,L:�`��\�IUZ1�,i�=ٓ�ز�8�&�Y�k��X�P��jkJN��Xn���5��ӗiq�~�b�wE?��!
q�9k���]�tw~��A`��u�X�1Z�ˌZD٣� �`ֿyO.�X^�����<�o+\�h��ŀ JA@bj=4�ewu�~�4Ʃ�,yY�R H<�@���ca��$c��Yp��˘N��߿��ߗ$+x�d��G��d��Z���(�Ƥ��>
	��#*L�_ٞ��?���ѐz�~TU?^��Fs]D�RV;5���S���5M�]��r�o�kK5_�s	��73�ei�I�61����U�d���J,2�4�,ࢉ����hre��_c����!����=86T\Sg	��>*���ְ8���M3�n�(T��된�º�4�Ô㧑��S;���,�)��B�O�IT�5�����,|�x�dT�+�(Y��UID�/^���0���X|��
�T�nB$/`�6������Y�Z�
��xe_]]���613��UF�`7�Q^�3U|�7�sz��W�r��!�8�v���yMMͣ�m����))���0��SN~���x��p�l�8���a�铱���T�K{�{f��FJ�r �)���I���T4���K0]u��m�(�j��!=q�0�	-�7�择t�S��F�L[s�'|J�W�Hق����@D���O�[��L��bm����(d�k�^0&��Z���:�0���O%j��A"k�b��>����B3�1.�̘T~�rHH�[_AE�~�V�����jFA�֋�Yl�忚u�1oZ�J�[v����0g\t�����h�K')�X@;� �xMN]ZT����'#q�c���C�i������^��b�|�O��>ӫ���W��y�����i�L���S3}{�$����4?y����߼ *ܱj�����q(D�@h�!����H��d�_����.�J����\P#P߲��WwЗk`E�:u�9�9?�ː��Y�[R�S����]L[ԑÄjƞ<�Α�:���ޯ
�q���W�b�o������A��Iu*�#����o�-��ӫ���:�ٶ����Ĩ����EY�МMEs^Of�qq^�s0u4�G���e��95l4
[;��H����h�o�c��'����c�XU"4VE�=�3.�����)LuVi��L���@� *Lٔ��#T˯*o��Q$�\��8���'wt���+� yrp25����hh��P����St�?���3*�k ��y���B�:Wj��/෉Luy���y��h&i-w���ыR�DZ��S��^��I
j���9�)%�sD�~N�ɴ��6�guB���]`M�)r�|��C���tdG���p���b�z:���EÍ�%��U��C������Q;P����句s ��EQH�h�}��~_=��L
�!�C�8��^3$"�a��^����z�^���Nuk�"MlG�v�������-���1�������HJ�צ~���}�%�F�zDv�p"��[���Ӹ�}[�z'$�Q�h[XAgL�!�"I��}���o3?!���)m&}���Ph3�w\uZ�-_"4<��S�����R%�J��}�����FgAX����ͨ��&A�������ít��;m*�Q��!u���������ު(Y���f(,�W���C,Al\�y��0�j�3�0)D�ܸ��R��������#&��R,��a�IC�ۑ��.��,|�NɪS$R��Α�6{�6�Wc���Է_�����:�:�H�x�)m:��������1BfVf�۾�1�[FFF��C����Hd?����Ȏ�04�$ Û���x���fk�q�ؤ�hxy=Ƈ4��t������E�r���i;��1c��w���� �(i�f�����Ld�*��f��9���j�n/��B�>�M��f���R�Z?9�F��y���)��kiii"��GZ#������SA8C)���'H@ք�z�:�#��'^��_d�m�z���͛#8%�����(�z�$0wi�G8[���\��U*�!~H�ؙ9vT�Պ�������(.v���āpän.�Tw!�d%A�h��\���"��hV�:��./#���5޵&�k=M��d��~ʜ��D�4-0�œ�!�3;[�0~�&=\k����^xԙ���rY�#V�r����޵�C+��'E�A?�.�O��$x~�k�p_{�p���c|��9SZz�߰x��r�,~G@�w��dN
�Gw����^��uAQ>�O$�&���+���]2�2t�?�� J��8�7�`0?1�$]��`QJ�h���!�i�z�/!_n{TU�p�z�~�(��%�;8������r�J3�C����kze����ճ�ee���{t��8_��E���ڲ��
����3ܮ��K���.Q����esO/%�����IY�|�U��!p���nԳ������n��|��r����;(��"O�|�r��u*L�V,�*�5�����{�M���s�e�N��Ze9
&-2y�[�� Ex�����q��W�G�З���W_c n ���]U��xa��څ�J�ֶ�>�88�U�>���;q�f�օ<p�26���3� ����·w[%��z/6�s\Pˁ�I��W���D�y�rVD�M�.P��k���s���vD�Ҫܵ6���;����	c`}������Ȍ�FC����͸����Ύ ��q��G���fq�2*nT�^0*�1S�MZ���������wu��4Jxc���v��w\R%�9f	�=��v_3��El��k��aDO&�^I_%��xH&��=3����ϧ7H5b�el3T�2m+�IM�ܶ�
�{�3����p��3�vA?��G|oZ�99����(�i��%�>流��3���t��	DQ�I��P�\P�Ɔ�[����G A��L2���{S[4BC�y�յ�5�=B��Fݦx @i����Y�68�-21W��1��6�Ϝͨ���:���h���i�5~�z��zp�0���	���V搗��$�b7��ɥ�ff��ꦗ�[Ue�r-nXLE($�qI
�}�!�na��K,&��e7�8�`�55���R8�������em_���g���7���[�kPHxg�?�\����#�x<�D��J�T�c]a�5�-B�$� (�t��&!R��ŏ1{�� 4 ��i�&��9k��f�����F9����a2��vR�h}�xN�� !����X��T���C�Y��k.���$ %SWS�Rb=s�º��^�C=U��j�>pv(=��`��A��B�ݏ&uK�1W�gh�,��k�%P�I���a ��ߞwQ��w�&J#��oV���w��7"��ݕ[+Q�ح�"�e��sq��.�4��;���m;-I�Qq4��n���T���WײΪ��Գ����]�`�4���b)���Y���A��g��C�/�֌m��X�>�=���?�70'�J�?D�ʽ	�t�a�@�aGH�=א�Ժ�*�_d���Y�@�I3mM262�U�7��B{D� (�񬓜a�p��݇�����A�\^��`4��txw7����:�O��WDL�1�4Ƽ�"��%�������S�E}���`k;��u>~3�Ln?)�'0�:�������Z�ёCHH�uG/���'<<I�
A-aN�d�b�j�'�E݈�������@�ni�6�		~���X�,s �u��`z��
A2Si����ݣ]��ăA�@��"++���{�7�<��r����
�y-/aX�I�j�c��L��.X�������V�
�$W�*AW�I�=�l��X���Cs��d��EשW�_Ys��'��M�cd-d�])73�g�� �[-�ʀg	8I�7�O+�Yz���-l�MKKR�ގ�ނa�pԇ�f�Jd��ź=��O��w����Z����3� 6��B��ݪۊQ�G��R��%�2{Dm?ی��ݐ0.ᄄ�#I0��"�A�2GQ,�l`|<!V@�D�.&�����>?�s�J�`�Cյ��������-���U�9e-G�Gl�R���B�с�R�|kG7Z��V�Y�&NMe6 {4��q�.yAm��|D�l�c(~�[�{����ڪ�5�D	�Q�AZ�7,�R4�I��������^g;e��&�f��V0��N�1ӵY$�y3�-K�B`�N��w�V�����P^u����įo�˝	���{�I$>1�
����� %����˩W���p��"��M��S��޲�j����0�r�.S#���z1�UVR�4Fz89�_�,@�ݟ�))>OU�U�;LT|�<H���0��^WJ��������ÃؿU, ����p��WN8Y�z��R��� �4tTC��[���LIE�n�B���n�eN�ӥ���?X̆��tf:�ܟ�P��� +�=�A��*+�M_嗿�q�R��C�G(+����D�2yJWQ���]t�N)�ڈ��僝�;�.�@Βg T��6��L��@����q�q��H*`���rrh ő�ï�N/�s��B}z߇�bAN�!��'zPn���Q��!ӧ)ɠy�Ig �����N�4���+A��y jr��Y�0��A��4v��5��s���~D������`1!���OgT ��E܏�U�;9�ܦ�v.U�ޔ��wR"�ޛ�_��Ａ���P�@�!z[��y�6ՙm1!��.�/Hm���s�A���*@�	����X��������u��|j����1A���K)��<h�5?i�����둔�Y��`Y�{���2����������;�1��w�q�=��ԅx�\��<�V�S��T���3aO�d�#�$X<�=#��U���!��b�$��-��Z��A�X���oK��҉��{R0�7y�������Awq[[�:���/�b �'�uU����&�$'�����o/�g�� �p�𐰊|��Ѻ,\w�� 
OC8��k�̚��©�3�Ԝj�|>����)��%��15d������P3�(�{rv�9y����?���&���a��r{{��8���'�R�]�����9T����8�5K1���QW�$�}Jbⅈ+zɅ`;�
Ђ��_��/м������v�����Q$�{���;�0�t����-(i�RU�%��iK3���C@X� ��@WTD�Z�F�H����EH�\��dmo?��v8������Kʨ`������\��{�a������Q�3_�I�!U���mbSW�-���}і3PR����������)OಟŶq-�q<�+�@)���/x��Nj��H�~�[�M<S04���"� ��b��>3_P�JN��w�AB�s��~q~w�5��e�-f`+=#S��h�ɸ�=�	�P�����")��D.��m�=D<w�O�����iz���t��>����=�jw�I�]�,e����_c�v�lv�~��~m��V0�DrT�=i�9�bf7�_�MX�g�uY�a�5��TE��Oٱ��6��Q<���;v�JaBGӓ�۩��.�HʹZ���#����z�8V�~��(���ل�
Ŗ�l	�=K1


��w���4g@|v���hj��`a`' ����K�}��u�1@\�"���B̏T��QU�I�+�^���U0(;����-�M�xbe�Jċ�W����sO[}X�����Y�y���$2}}�v�Ƈ"��=6��ݑ�t���k1iEz��MMi�0�8Ziz����>0Y0����j֠�n�3�"�$��f��hg�� &�5��k1avZ�7SGُt�x�x|�_?�H�wlu��{''��ko�_$��>��>�9��1��_�]��&��p�d2�DR*�p�|	uu��zүJ>D�q~^vttԥ���:!($�l'�:?nAJ�EEDb�我_h�Et &ق��NEGG�GI��^���7 ���2u���7d4�������=�P�=�����X^l���:�u�a�͐�tr�w��� m1�a�m�1�/,m#��k�|q�^����	%��~T܆�R�c��dw[��uj�u`n(x�.[�/w��yC߿/��V36�|`qQof���)H_K��$�v��6�RSh��펿S���B-��k��'�S:l��K�g���h+�ӿ���(��7���������i�i;�쑠��%�a��zf_�gQ��[�OW�onOG��ġ>��=����3~����
�{�Ȳy�g��y���{@�\�v��$.�x�2gML�Bsf)�xǡ��=�'��O��w	Hu����z�-%�\wS �%tJ#5xzMO�WYHѱO-�tj��������}�+�uFk�K��J��ʹ�p��'Q
��R��8)�'����>πt��2� �wk�t���3ҭ����"�p2=��B&��0��3�Ԯ1��㰄���R�#\�!z�v[}��Nw�������?R����s`b�U0N�1	�̛���+A
���Q�5��n�3��jc�������Seɏ��$�{�>pU�rlzn�VQ[�=��ly-�W���GP���r-����V�ևX@�	���a-Cb;y� ����^V�����O��=ҧ:�S�~�s��E�p�������i��V����o�r�ռ��fV�@������D�t=�7�����\�9���D�z��W�]A����x�߼y#�VOedJ"@pܾ�9F#[t��*g&ޔXh�D��ĸ���w�Ӻ_���͠����_�1������>G�����v��LIy9`�����#:50��h���gY$��$'�^ �\n;�*���_�|�GG*�[>W�q޼�0 O `o�	��a�F�Ccw�4*ɯמ�7H���k�ӎ���\��]U��m�!g�J#k%&��z�؏F'��e���Ot���4zd%����a��[1�K��K�4��?�����+s�T�,�VW����|K�H9��V-,�Z�/�4�y�`�XB��*�М�H�XB:�$��}ڧ�">�ǻ+{pNY[c#��?�J�,�0��Xr���t�@.Ri.��V�C׶�*��?T7�%z����(c 	����N����"�T��t^�M��nݵl*�][����U"柞���.e��\����(%4�'�}�����i��Ů���d'|� �:=�c?���;�)��,(~���:ҷ;V���3�rp4�r4R�}�è�������e��l��_�����<Ȁ���+���KV3s��I����N�_��mQm������qŕ^�z;3/ Q�e6��_�/o�����F�_����=[���O_ӎF�k��z��q��� �7ˌH_fN&��1�U=�2����A���v��^��5�ː�����nFFFd��V��@"\�.د�!R��|��mw�@� r�7K�?ܮ6���^��I�v[�ӎ� *R�Y���j(�֖EH����6:�*�H�� �`������D$�Qx>S�9m4�	�kG�ҽ �q��ϐ茨�B��R?�a�ZT���b �V�5c>%�mC��5ݚ�l�����z����(�kR��vtXө&G�����O�^9hLYE�� ��i����k _�}��|�&zz(J�o3���5	s�3�0#L�3uW+C�u@I9Q`*l�|�Jo|��9��>^W��ʆ�BpDEEu���q�ă'�'&�0��3�˵��=�}���XW;�OlIRɂ�檠���m���ffc)�Z�m���Faj9�&6� ��g��=�zDpi�p�y�e��{L9q����l�m}�'��À��{�Rg(���Z, �s�_�����T��L����ݡә+t�C�������<  ��AAE�7h�-T��5�%҂+<Y�E���J��Wz��9S�pss��f��-����������|Ye��&;C!���b�V֘�7�>� }z�w���CB��8<���.��9�w>���YY�9�}Y������X[�襑	5v���T���ʍֶV�o]�T*w�y3�!x�E�m����DJ���x�f�A��و�)M�=��zR���I4��&�*Ԩ���=�O��Hz?*Ӡ#�ME��\�JT��)�oOo��N9�*~G}���XB>h��Yc��՝ꗌ���77��_�k�`��!�Βm���L*����6d�Xf�Yif�.�*:[4��*2�!캍>cˇ�=7�ԟ�F����k��^��݊�*d:�Y��dK�S�o_jw��ckw,K��ȳU��F�4[�C/ ��M�㋆���R���Z+	��+�f����3�����s�\��O��!�ظ���!)'9�Sa�0j�ΨF�V_��
�c����8=.�[�|u�୭B����}/�W/��5�NG�r~r��#!�~Θ���Ƙ���w 	P�{�<x�ynG/��Z"_�k�����@<LVl����00����A#�tMuxxX��d|��3r����iS��Z}�)�=C���n�5�	����s������Fp����Z�BK�گ2�B�u���K�8�m��_��)v&�:�Lu�[�zh�n]�\��{�c�eH�v���V���.�N�w��ͩ�u�ux9~�e��fVX��w� ��5�}���#���fʔ/�d/ߠ%�_H��B���?�"9P�k���]�m:��I5[�n!Y19����Wi���F�ͨ:DE����WԄE�`�"$�89|��~��[E,r�KHVA�1����-��sarv1�c�vø�<�����O~w���T�������6
�rF��̺`�Tw�[�8Zhw�TY��񲵃Cؘ����{�N~���"�Bu���vx�I����|kkKWWW"��ũ�F&|$��⺭��W�7���ޕZ��iG����a�Z�[<�vɹ���{�M��c���>]QY
H6��mI��7H?Л��p���w��q�����ْ1Q4����&K��ݠI0W�r]����!J��U=q����5�����8C��' �˝��_~+p���Ė��G�<'%Ƽi��~o57�t����tj7Ks9�'#6+��y����m���8�����((`L?�aɆ#���3�鲍�%k�� ���X��i�L����8�B!���S��%���E���<�#w�!��imqX�����)S�~}�ձ.-'�d��q0�֔��<?����BON�Ȱ�[��5Oi	,��¶�e1�uG����0���Z(?���l�����/�ɾaH>.��{k7��J�u%h 쀠@'��#Zu¬|�xX�#���B�f�3L��~����ш%����z�7^R�zg|����נ$$�gm� ���}��%��eJ!QZO��w+��P������}i�X#E#E<�>��Vd�C7�M�*.�k)�}���6�L�Q+�+�vX@XϪ��_��d�0� l1��`���y���{Qm�6��?*ǀ!�Ӓ�l�3�H|��e�}K�~y��nggg��b�)c�E����X{�1� xV'l�E� �j̑LT�� �T�=��(,,Tc�fk������R��*�Q8��%Y&�ĤP�����F�8���m�����x���|8 ?�(q�n}����q#`P�V�3�QԆ�Y5�&n{wrr�s>�Zk%]��q	(���*�W16>�X�8.�,9%�|��s�EiII�LE�To��]��b��=	��<�)����w>��w}��D������'	ӸO4�3`K�α�������?�lw����ׯ����ǔ4�]�qE��8�����<���Hd�d�fP zE�,�@�O���n�j�;�7���}E����L�}��O�F�DN4�%q�� 8�B �� �&��1�]hM����w��Mt�H������GX*�埅�g�����{D[�_�퓏c'� y�#p��(�l��(�r�X�J%�I�Q�� �t��?3̙{A�����8�a���]�����z�}^DO=+Goy@�ӊ �nU�ت[>�jED@v���x��8e��a����j3-��hݻ;T�
��1���c%�ԯ4Ӎ,��m_c�;C&[�o�麲��f��}��)mT�h/_Ɩ��XQ������H������5zqc�`��N������N���A���6Po=�}��$�!*�H!��=I��X���9ćz����8�,׻�OlB�������$�)a�r��F6�y��J��l����0��tv�C��B^�	�2+Xffg�aN6��G-���5�-o�6�$`hi˱I�����յ��B0��y�R��������uUa���^"8I���s���O���A������L��3�����]��~|㍷��n;�����"����밂�g�|<��>��_�jt�,eI@ߛ�k/^z����{��j�Z1���G9�Xy�*����k��s��-�= 0��>))���,�W��9+#���I�R�NYII�6�^�Ό;ֈ��-<�9�H"zb���S���N�����]2��Q#C�?��ѫu�4��8'��'Z��x�w���x��;�e�Sd,���Wp��(n�T�.����	.� z
��:�!7��?���[O�7h�1��)O�~�0�wx-�"X~A@w�@=h� ���=惃��!���K�6S������h��y0��L�o��P$/���=�BA�׃�vv	YY#;��/��C��i���E	���;����n�'5�Sy?��dhaD�~�IL���I0�Xf�Z�ś��>gE�����/k�V�- �
���ײ��`�.ڂ�@�XX
�=0�q�DR�r�L���q��a��}��ʰf�{�^��Wx`b�)K���~�t���>m�,f��h����)�-L����R,]%Xf�h�Jy����^��*�d䦀<�A����n����T-���$u�Mp����\Չ}�=���G�h��=�&٘�-R@٬�|"���k����Ù���7$�H�TPnV�{ˏor|��I"�#��s߼@L�������Rd�~J��%�Z~?A���D���m��M���~wQ:KKG��2ꭢ�ӳ���=��Ӳ��݌���b�'�,���� �Se���g(g?˪[_�۝�
m�-�I�Q�.(�+q�/������!N��L�b�!�U�C�M�g^O� &^a�s�o�4h�xث}�8X����#*A)������N�skH�6�֯.���nq�h��#T[�$M׽;Vk�#��3w|ƒ�J��^RR�U�8�
�?>�����Бdi��F:���'��ˣ�B]VȨE�x�-|�ݛ���1��xsQY{6Ą�5�s��2
&0�v���J3I��Q?7�)#�ZmP��	??w9
�6�L^J����'^\V�h3.A��湵��L�$B1��]��a���0C}��q�M¡���\#�w��>p��w����3>U���-M�9C����g��&��*>b;G+��psK���Ք����CH�K�x&���ˢ����[�-tX�nj5�W.)�6��<�a� }Xh<�(O7����i���v�����+l3�	�H`*��D�2��%D�t��d������]܀��=�1=��fXXY''�d�&�$�Wq�ޗU������������j�+7 ���X�c��+��������+ud�o�s9�0W��!���?˥�&}@{�3�+}���jG�ɘ�3���S�crJJ~i��,�osb 	 )��Ӻl������H^Z�an�12�D���-�FϺIc^����`�nԠ����#=��K.o\��!�#8<}#��ƮXc�&�l�do���h)���Ψ8����YsI33�V_����F��^3MNL-e��A�{��������cR|�����e��}W�QB�Wh=yu����ٿ�7��MJFEl�5�<�C?��o�����U�Hp]�Ԍ�wW<72y���qJ&�������fbr�ծ蠑��`�Z��]H	�O�H���Q�AkM�^H&��㔰rGc!3k�{��΁�*��q��*��/}�[�{���,A�Ү���jZ���{����e�Q�ݰ�>�4���OP�����ǔ�7���!���PM����s4�
,=�i���a~��z3�s�-�����3�lQ�j�OUXV�R0�M��$��u[ '��DV7�A�a��NcE/b'-���������g��\)S��m>6p���������ظ�<v�ᴨ$�/Y�Y��0��"�����4�T%�����"1������¡ Ug�[d��vTi�^��ˇyZ�֑�����>^�ak���>�6�,s�����ߪٚP!v�HA܄�E_{��K^r�G��H�mo`�
~<n�Q�y�`�_QJNN�Dӡ�*$B	�{�����;>0Irwfe�C&7���^N����`����
$�v��Y�l$aaa�5��	��WEW��0cq���Tx^�}0ڴ��O�-om ro;�Kn����$G=EE��6{����weҞ	�_z���/FEU�`��,��������� <1x�H��b�h'���y��gcӞ�t�a��ݎ-�?f��p��L�k��PӦ�d�>j�7+�ҚAsay3����T����M�v��	*U��J;z3����Tc�c^V�%E \TnA�HV���о�7b-��}�9!93?�y����LGQ�#mk/�02����������%�D��xN?d�ȉ�bJXX����t���o΁Hс@�zb�r�v7u��%�5Hה�`��궾��}�g\�����Zw3* Dy���i I���RHij�<
���i�yo"��9(�h`���p`3T����-���*~g0܉��Q�0}E���dgg��~�v
����ױ��vM^���Jz�D=5�m�w��1 
�$Ml-{����~mc�]-M��w��뼀&$��-C�V.��w��}an*�RŻ��u�6��/�N�A��ԘV�S��|�N��YU���7˖�gi�G;���Q(�B4��C��N��Ųʺ?t�[Z<딄M�{�ۆ��:�����ܒ�L��x����d)3n��p�G RPM-H�8P�g��<��-r�LFǞ*%M�z>�y�v�X,`��S2�D�!�]~�mm���}tx���/ឲ�X�סA��֨L#�G��j,�EצK�2��|X����o��x��Q�@N�"�����B�'%�6s|��4~ �8Cp�o��y��)���)t�zyl�,b�����+7�eT�1�J�4�r����G�[���f�Ԕ�]Y]n@��JN�h�FT��_d	''��If��5�Q%��o�m=��������~_������ٟi6�6�R��j\���L�^��Ϻ=�e*++�z0q��4�e��'Y7?7��H?7���P����l��bz�*r�K0E;�ה;;E�WW�D8;i� !AVTv�:�[x��i$�W� �c7���=.��i�W���O�\�|���]%�Z�K36/m:]�e�)?�F��,/#���-Y��i���y_�:�UHi��enL�~��C���B��*�S������an�m���`n11Fk(����������hxx8��G�A�TT�'����@CѦ���0��vɝ�����,p�<p��;:^ +��ܟ�n�}������ĵ���@I|�yO4'����T����_,��65Ɖ�z��ϑpI���1�bpM�#��Z��uP�"AG��Z�kR�j�2e���?զeL��Ï�)'�ӫ���l�P���M����י<�&��(p���勣.���bCw �W*�X1
�w��o�el��Œɨ�D��i)p
��R�)����~��5�jPQPl����c����y�X����E�)^5�P+F������%!D^�Sȡ]��*Ltl���C�9�4����yM�����a@�sC&�ĳ��UWWn�K���c�M2�����CJf��<�lW�c���#�S��?�]:�%��6��c���X<�qK��cZ��_:킧��ߝ%��IHҞ�rw�R�U,���3`�E�Y8���^�@��y��}!9��a~�'�?�R��r�L��>Y��J�#h�I������{jl�x~�����W����T����:

�׶{v��h,�r������p�cl��sZ�7�ڱ�ѽF�H�-A)����W��y��av��].L�͘�897�o��x�: n���6
��^1���"��"�'*�ə�f ����Ϋnzid����\�w�\���X1I�R0��U�C�{�)�j�D���(6��N�q�,AO������vK�wT��e��0�LW�Ha�H�����OW$sR���m��ݾ������Y=����O-����[���q�*w���"0-n��_���W�$1����hR.�}չ�ZG�<�S���*�'�i8@����`î�.�s'D ��T$��ta�ȍ�	�i��Ѩ��:-)��@\�~��G���㰁�`����aŅ]f0�$D��}E��W;:��v��C,Y������E�3��b��Y���ϼD���~)17i%q��qg��h����V���HO�
��联��X#g�̣��G[��˔��~e��JKF9>�,ZK9Q�'���1���*r9 \ǀ����+nw�p�B|{��3��(�*�?��q�
f4�[��YK�}5�����1���l����?��v�&O0kC�8JTƗ�
 ��q��44�+ʕ���u��W�����֑eѲ���H����8'�ũ_�~���j���:�(㣶�m�5�|D�Z�$W4D�wR���ȿ/��z���7�:R.$'�j�߆�?�iH����.���f�Y�N�u�����]���g9�4��,�� ��\���O����+���zΧ���/���o�Wz�#�Q&��ʔ�N�v��f�v���	���H։ʈmC�*��W\���0=�<�i�ZM]oh���k����_���)��1m:,c���r��(F��C%y��l�b��C� z�)�D�dO�c�n���<Bnxr�ԄU�^^�a,|��瀩p"�ŝ"̆�%����3������̙����()��g�ι�OL����⧞9�w�P�$�2����P��[A�DO���D��i~"�q���xp��ł������t6�
�I3�)��"9v�B��h�J��\��Y�����/|:~Z0�3޴�T��*�������2�'��4}uXT��5��J�HJww��!!Cw�H� 0tw��C
�{��}�ß�{⮳�Z{�ާ��$]x]�ʟ��H�(���*�J�4��F���.��.��y�~M<'���}(���l�k�����]pj�:>�����)gi҄�S�X��������2�0���Hmf��K%�:=���ocxt{p��3�Ĥ$@�b���ʦ�ͫ���u��%`
5���A:�%|N�F�@Ԋ}g����o��/O�O�Mp��������g�� !a�i���yg`���\����&��b�Y/���a7�7Ј͔�f�e|��_!����|�h8P��4ɸ6&����/03�TF~����V�C9�a��[66���֓�x41��[Q(�IЇ��E`���^��i���t�.A}�y�&ɧ�� ^*$C�8a>f$��G����מ�'i���"&%�>����,����T��ٖ-}u|� �ڢ0��]d+V�%��TCA=@C��Zp����[X%�'������O�v�W7�"�k1�y��ןx�y�j��ޟ)ji�t��F��8995َQ
�}~!I��?�	)m���LRR�Y�~�(_�KzC_|����7�w%��
2TX����))^�e�esXm��{z��j�����#�O����D���e �"�cv�E]�hy���U�#����N��ڤ4Qm�k��3��qS��1�ׄ�p#���Ζ��CrK� `�s�syh��65Sz�����M�t��|��ҟ��=�t��',��|�U����f׫�1}��{yF��BXH���� �3a�Z��p0�-xf:�H:::5-���2��3P�Y�}�l7V�Y�X
�y0��%���
�
f���S��2�nP���*1r��t����ح��)ߗ����%C��>���D�)�_��f�6�fT���"�F$�/%Er��9�V�A�8�s?A��>��ݥ��d20�)��^�D�^�Ju�/���~��^���_U�*[R�������a̜�=֞Rg���%lpȢY?#*�iK�V/�ˏ�^}����#LF��(DN��L�8��f%(K�"��b���r�T#dR��a�s6qM�J��Y�G�v;Ƞ�jTQ�P�Rf!����[G9g&�Q� � D��מ*��zu|�D�#f=�G�J��iCrV�zI��t;/�]E��2����?vȪr�<�H�C��A�����0��n-����&�[d"�|MD,���ͩX&,��nR�ȵ0�x�N�D_O���'?Y{�͝���� O�j����6~~YYWc�ސi�N���U�����A�����ce�*1-9��@�p��~O4�否�����{w�Gz��|p���P��"�׌���y�~��Sg_���1�]���F��w���*T]]_�s�3�L��'��z2�G�DE�3S��٣��]��i(,��FQ]\��MP�h��椬=���	E���GC��^��@��	#43�F�K��-�K1����q֘K�'"�����ATJ�MM��� ÿ���%�C�X�.��5�y������h:��&�gj`,HOˇ)����Gj�S
���u����Q�A��VL�h�A����0��/}db�z~⻲>�gp��H��ރ�GG����������X3#�2UX�����lO�mȅ0Y�P����E%���Ģ����l����gh�ǚ��*{"x�ᅼ[���>�[2ݙ�������tl��$��u@���:՚���{��l��b���/|j�7J��[
�?v�P:Za��?ݗ����
�rL�>>��q-���O�̚E1[T��0șwz��Ł�	�z�a�ؖR'�ݴl�|�Ϫ�Z��dp�}["��y��zQޙ�����%���"������|R�1�̶3��VL��'�z�����-�x4����k����8���C���F:/64��H���{@M+k+�t8�k/[�����.�G�D�:J@&�Z[�ި?�A�C�_e�{A�XYY+kꆦ�VK��Ow[��Z���U:��X���0�\��tjZ�\�a+<$c�	���|�@;��::��.U��(�ww�.4�� ۧ��C�Αg��;tnz���f�V)}J �ӗ]"�� �`֙K�+������s�A�����
�����BBr+E�U�)5��!��f#7g>�D��YU9�K������_�I???O���w�?���J�‥���K�ʑ����B!�K5��w�����!����|6{���Ն�&_Tx8��U���ˏJQ���''��p-�R@��T�K.zf�22��X����pf�J�pvG����|M����������+ �%��5���'> �7du�-:�z������}�L�,?N�2�N����h����/�-��g�?�5� �(&�)S]����83�Mc��|"��]�ʾ���DE�����r�������Ӎ��~��z�xM;�L;}��a)�F/���O�M��ϵ��~8:zq�b�L������R	��x���?{��<�Y�����f�L'�s �Aʟ��KD��Sb������J�%��]Z�]/��i���Ddx�([.�s��8����e�L/���3ns*�L�T)XQ�"�X������(�iN߆��ps��D�]6/�Se��5��������EO�Y �.�#Ђ�вm���y��k��x���_D�^NLt9���-�'X+{��O~ֈcG��SZff��9�xj��qvJ�E�/��k�GQ��Q�=)F>�
z�����쓜^���-)$*.�%��q�A=�RMCF��Oh^�0�eK@�M����m�����;�l��@���1L���ߴ�O�։��,���'H�B����W�k*�0�G��R��wX��>�� �4Ӻi_iVf���o[�BM���ҼZxI�LizY]���ӆws3dE�W����t���M�LP�[�)7[ߪ��� �(�������`-쮳s�zf�hKDR=���w�����o@)䤻m{�\��v�S����p�}�Y*`<�a���OWٿ`�͌p�ݷl�����R�߫uo.�`7g�1���#�Y{c�g��0����Q���Ky��*H &Y�������/�_�)�.&u�P".c�A�FVWW7�M����s���_YקP���)iyix3ͬ��g��$j웲���Oa�
���2>������HX�{Pz|�p0�b[<�|wtKFօ#�R��e�YX��[��ǫ�gP�!D������l��T6vv���\�>�#i�桁A��Es��ٳ�8��g!�H�~�ۼ� #D0N--E�׫mkf(�_k��*z���|��{owTG��2Y��D	��?��`�`�AS�H8�� ��~�XܶK�A�����?���#F�
��G͜�y�̘��_��o����!�U���Cz?vV����������x'r��7T�|���Q#>!��$Է_�݊_��p����'5$��FF?Η#����D ���RJ�u���F�_7D�L�\�U�����(g�������G��v��%�ji�c~Gku��(�����T힂@�ʪ���F~I��Ӻ���Zw{)�MC �?毭*o��8���C�����;��ި!<�.=�Q W-QyrtT�Ք@��`4���B'��Zl�4@��y"J�<��6|��4>���p�-/�E�v�S2��z���5
�� 2�PB�������CT|첽{:��jb�Go�d���v^���*���KU����t�#B�O<�� 33z�3=mq`�\W[�Xt<+��Q��cak9�Yw8�z�k;�����s��^�����jf�����mp�������I�`Nww�2U�Peu����7����'χ�y�ٕ�;���9�r�('��+QHW��e?q�yG�[1y���n���!`�����I��;�dZ"uk��M
�ҷ~���z��cIHl0�UȽ#M��la�~̈́n�É1�&��V��A�$ uY3��є?a���wԌ�$�����K�aM���k�Z�����,̡;fZ[3��	�&ħU��q���梍�Tٵ22�<�k;�H���y�mnNccc�̌M��Ã8��Y���|)�CG�
���yћvO�A�<AZ�©7_�{ry���[d�=^6ب�m�Q$���\L�z\��ot�E;	Z]����m_�F[Ѐ�:ӻ������u�jG�H�|}�!H�|�iq�i��o��x�Y5�g;�2mS)���"��JzՔ�2��3�Ͼ����_֔IH������;M���f��'g���C�Z�����{����R峓��Q9�`��������T�?>��
���_�0B.���^`oX+��������0�"�����.�`���I�X����S#��t8 ��WV"49������:@����teee81�\ֳ����5�	C�����vWj�RTe��|�W����,��b��O3�03���g6��"���Ev/,�]�^ �Ϯ�)f���4�[��[����S��BG�Cg�,������A���Y�(�H����o���X=��?�_ȂϢ�n���g��wʡ�>��q�㬭G�v^{���k�ԕ��ͮ7�O�u�1��[[�{������t�ī�B�������7��ȑfpp\% 
�krȨ�_�e�7U��!�1�s<%cO�������"��w���t�.g������<��JUN���]�J;��4sri��	#���џ�08�D�-j�IY��|�.�R�����K��cHR����1O~��g����T�Ľ<rሏ��+����t���.�߀������4�@����(ڔ�s��i)TLT�p�~<φ�#�r,��%V��v��a�u�j��]Y�C@��g�pƳ���3ۨ��+���ls�*A!A���;������J�˗�Բ�o ��"DK)�x�<�-���D�s��}LUUdc3EY+�Y����(®q�W��n�Y�;��l��#��W�]&�惹�/���{��R���G,���jrDi�EA�]O�D���b $8�m�r.��a�e�4c��DEi��^2��!�R0�������V��Ih"��y����� <�c̳��_��?���ڿ~�N?�鴜:��͕l�F�y��M>'�M,�O,��x�6�
=��~��Η}���o�UW��[4	J�p��W1<��C�紌B#��LG@S�;(�K���v
£�p���A� )��)-혈pg�)>��!gxn�<@��,l��bZ��b?/��@#@>����us�φ�Z`�y�ͮO��_��6�1�����7/��k���\�Z��Fc��Y��{���
��MG'��\���)fNz��kOXß�	d�[�2�(]�',��vò�������c�3n���E�|7�9^���L򎗌�D�������G��]OL�l$�h��Lc��\���7�bץ���^�a���H���qn��L�2��x�.�[�[�_�%�uz��~E���ѧ�?�|}�	�V�w��(�2�4��?p�w���5:����wjii�,�p�@��ӣ���6t1��{Y�ݹ�pymX����Y�.P���r|N���7V�+��X�׆�1MzC�u'���e��Ƿ=
��P5��~#~�6��`�m�n��)��L����'I�Y/�e�����$���[��ߟ#{�৴ze���);�s^n�;m'P�
JD@��r�w���S�J��Ͽ�i�H��ٝ����J�ߋ�ߏ�#t����fdf>畒*a7�ӳ�oumG�.�"&���f�Z��rrrlN)�j�9?�N�̐��֕�O�#�k�o�h��\��K��T��:��6Cb����v���i��{s丸��=�M�Ӊgd�]����h�&�����q{I���c��hnN^���˶�h}����8pJr2#c3��I�{n��Q��+��nv�|�.JS��H��z��N��)�x�Q�;�+c1�^������L�PM�H�L���s�$�F�1_�k��]�.<8F�9Z({eh��9�W�*ӄ�'3+��<����cs������E+|x巷���zRR�ܨc��ŝd�^3�;٥ؘ��]�oB���qr@���ΣW5��ߞ��ٿOV��+���Iz��Q&Υ%b	�����DQug&����%5e����C�-��$o�ԟ�S�c	[��4����j3��BzJE������LNL0����"��Lg�H�8��к�qr���ㄮ�����N�43�FCtuA�3*7; ��::�%�\��ngٲCB�1�0�N�Eȇo��u?_�H`�����}�y®8�@i��Ͱ��]o���j���
���+I�q�N��K��E_�=�T�3`����K^1��i�|#	X���3�h^�����/�BB������Qe���y���n���X|���a��2_T��;h$��I1i�o�UԂ �U���2ӧX��E�s1���/�^+/g�o#t�(0���)\P>�^K�ͽ����K�������ļ���,�1n�nж�pQ�S��Mqھ��*FrK2����l��>2Wq�%Y	��gga�t�\��oMz}��GU���������?.��rO�0�2jG�k�C�yJ4U�K�>p~H�eO��2�uSC��`��7�l^�����yll��������#$��L�,����ݎᣌ_Y����Q|�cc���ǒ��?,��f�疴&���z8����ɢ�� �M5���+��5bᴣC��J�pf(����E����G{��M����%i�T=y�ⲏ�di�V��Z��i��Q��Δ$\�#/䕋Q6�q_~{����=ӆF�W,0��,g�I!w{d��>�\\��ܤ���W7}�֝�_"rs,�?�ht��7,&��D�����a��R�&��ݭz���C+Tf�%�u�x{YZ;�Ma�m���"�/Jo./�,-雛��D�m�6��=D08_����C��YH������ޥݡ��O���1�_]o0������,VCJ"r��Cs3+ ʉW���2V��o��ɍ_�ɴ�{h*gE"&%���M���F��jXfhii��'�dہ�l�{RD��!�,'ʼ#�}����>��E���~�5:�K.灳��uƭ8�+���_'�W�8�	�U�^��q��T�!ݯ��GE�"Uy���4Z�*�;�J�h��w�L�U2�P �c�_���`�������x�!SC]��p��S.7�c�ԗ��aťr�I��O�	D�:n��R�WG���3��Օ�/�j_�q����5o��#,�ګ�M1������J"��ǭ�V��Wjt�l�c�"��:�SEaz�����$a��ڊ��&y�ݻ?o_O�Ц�Aݺ۔�G���'�.,��а\����G����������2	�C�4vs����Q��+�w�|,�_D �uA��C �dOW�' "�p���TbK_򜔐��k*Q���و;"�X�M���K=��������P�����C�B�6�[[B=��ɷ�Q��жֻ=�4��u6�M���8Ώ.�a�>��;s�)�����g�羳��(XJ�H�ܫ��"�pw�G��b��-�y��+��m>"��;�����F ��f�;���#�7��f߸���� ���ш����;ߞ���G�::*S°��ί͋���� ��I����$pB�H��=�WTc|V�a��V��y:�*�qw/�9���?2�hg�ʜ�z�'�=jw�)
J�Kk��w�=Βn����\ l���������(��F0g�n׺~"��QA�b� �|m~�b�p�KX}nH�A%6�Pa�`L��&�b�vʴ=f �s��d袙t0O��-�C��_����a�I�%��W���I�"�#NM�)��*�U�2�:�1�^f�_ʆe��4�>��I��]�F�K��t���xc.^��%�L�9t��q2���_�,c��/� ��Zgf|8�Y�|���� ,���ɒ��d�u�y����󀱑�nw��1�O%D2&�������`�����G?=^l��1W�}Cy�/�
�f�i�G�mk�P�ay9�O<�3�0	��ؕ0�˝����~q��,E�K�^ka�\�w7��`�R;Q���d��b��v��Ub禕R�L��v�\��0!_�tjv�9����nP�bmk	8�a?�g4�# P'����̝KW�T0t|!��5��z�M�#��  c��x.�qۏ���C�~��˟�N��c����x�򿖈��0����L��Ǻ���4�2v>��3��P\�B1*G
n���Ӧ�?Tfff9� 55���;o���a��Ð�%��ի����G�9Y��B��!���H��pvt�G;�B2A��>��� ��x�bX��z�Yw£�#5]t��P��1�V{�U��BfV@G�Gz�vZ9,_�9U�Q�Jߩ=��B53Թ"L��rf&���#��e&��_���',1�X����\wC����&"��8�E���lÏ���*�� ��K��rLF8���ĺ��ח|pHdN�ĵ��yY6$H���O����I���>�`�L�JU�ʰqk1JB�k��dD����|;M��߮�G+	0����-P"�D�� ��8xx���C�	GԦ��wP�Ԯ"7���@�[�b�t��m���-'�zA��`$���Z����¥����EG�E܄Ž����SD@�[��[��Kt��� (�r!�|�^ ���{��S:ߎI��n�W*��}��I������Q�(���]�ɞk*��<ץ��v���UU/�D�R�)����s6>�����M�������Y�9��{&\H�#r��$)��ζ�h%!͞�k��g��xj��s�@����*�nn���V�4��b�o��.��WV1i;�Nw�v4��������0�T~��M��N�h{"ꚪH������_���m=0<Z�h�>a���Α��2[������Ē��u4�J���mE�� ($��O[�r�Z�Hm�$��Se�i�<�P%���Vp�U�v���o\6Vam�=�\T4}��I��i{t���q�h�@���I��p{z/�2����ż�yy��9�9P0�U����p��q��nжd�yН��|�w@x�YQ'*�#?�f��0���Mӱ^��-�����疧�]Ǧ�%�W��DQhh/l�1խ�V����ɐ��QE���3AQ}+%
E����`�y�M���͛���Ð�vρ�����7�I{������
�����q����u����n�<��3'��Z}��IDLR�D (M�!��b��}�DC��lR6@^S%^�<��B���� �bx���o� �R�*A�I�M�57O���MC����p��a���l�W�311Z��2�>�}`I!���۔�0�H����]N�ƻI$9����!�6v$�kK����z]�_�0���w�3555���̎ T� <<\:�@��/)�����bT�R�h ��/"|�ܦc���J�hR9��8T_�J��)�v;p����s^.����d$� ?7;��:-[L�6�9v� �V#�<%�dy���42:�6 �;��c
/*zn�ɥ�&4�{!ݰ�a^�b~��bP���>��96H[���H�in�ʫ�4��"8�m�77oŖ�r�ebU	��0Ce�R�2��`4Iή�<.� �<B�%S�����K�,�+�/;����+-���|qZm���
g*1=${��Tu)�������J?zȡ�åQr�	N�=y���^��+�����A��4uwD�YL:��c�� ��Ύ�ϫl9:�>
9%���5#9�+�9ir�Gb(Zޥg�R�߭���(W�΅��[628���Ex��3��������.3$I�׹i麙���BN������o]R��2�ͧ��dk�6y���&T�����~F'�J�����SL:� =.�t��5�4�E=������_�us��a���R[��k�oWmDR�qX��H�.��j^,�0���3�!��������v�^�N��5úͦ^��ޯ��P����_*DZ���4�B�'�=�˿�e�V �e[x�������߱Ҷ!ȑ�5_��p��~�)L$?+r���:p�=0�oβ� )��;���^�U�a*j.AD�IBne 6B5m��_�')��o��Wv�}Dtq����9H��8<n����]ākv���X��N�	�=�]�	T��[�*�>vX�R�3a�7�$�$�R�O�����n%T�¦�9�7G��w�\&h�ET��|�R���Jj���ң��E,|�-�(~���>��u��9�a���ո� (@�3��l�'_f:n�������0�i_�Ц�����	A�P�:gg�8���c]}�����K���	�!�'//�kev枍M}�i�X^͕  0`ۧs��65~u�����'M�Q�;�N�����3ikkfJ*J�ޭ��6ݵB���%ߋ����k��:OE�U|4E�S��\Z�M���c��ᑑ���<�ֺu��aƧ���NڏJ���V��lt��~`�Tmaͬ���[�aҢ�׫y�D�q�o��Q�?YY��\]aX��	��&�J*��%���klrlj�J	}`������w��{�*����quv?S��I3��b�vjz�907��f+�CPj`�=�\VƓ�1&aމ�r��S�S���4SV$� ������!�I���	EȌ.��,(H�A�Ƥ͵{��23C�u�(19�r_��
lcuP��4���"�k��$Z�-����R�ff�X�NN�=J[}�����w<1��7{\sm��)#'�oHI�v&4_�^���@s�������2��p�\�����)� li��q���|*o*�=�+�0�v��ps(^��EN�jU�y����
�r��#)A�>�Ǌk���i�$S�g����r�=f;��w���e�3y�r7��8��\�VVŢ^Q�y��0R�C��8���H�z ��͕u$�I�Ȉ�9f	�X������4�.HcҔ9ܻI����/������R
����Br��T���F�����f�z�_���=ː'�F�J�@��W�Z��I��uN��M������RɳlŐɷ��_��TN~-7�3A�M�ɁwUw�PPPT��[XX�ĕ��o���0KI1������d��7Na���M*qĒ�rϮQ\(]�n�qd5��M9(����΢!�\�s=;Y(|����Q%��
d��.���ko���zYk{c,BGNA10�/����e���wpwW��~��x�u��'d݊W��B�[�����E�-��	��ұ�q�b���J��۟ʏ�<\���)�� n
8
L{�A�W�.퓂��?^��o�>K�dsu.��?�qr�줞���9�ɧ���rC��h�wD�%	����^x3��Ca�5sJ_��ۧ���i>};EN�'�|/u#���?f�;�f��,�y��J������5����O4/��4�yCU�2
��������5 �3񤣕,�S�K� w�޽{*q�d������^=~����(`���b��Í�8Eܟ��g>�$�r{�o��D��Rd�h1b]�9:P?ȏ]1�zz������5�����0,�e?U�a��#��	<J~v�e���v��|�&�B��u�Lv&B�[��dPD������;C0- <]���Пy�_�َ�(<���q&�F [��rs��z�ՑޟS���r_�$��w�%-�~���v���X[�-��  x�+�CȥJ=���J���>lc�������ibn$Z�4��7��CB����6�K���\~g��������e�,� )���3PQ;M�̈�玈l81�^����>�R���5*������F���C�P����VgXzϗ�|��Ѹ':��2ݿ�MTΑs<�S��t^$�p	낋���������2߷���}Td��w0�$�rrs���R<ڼ����'���ٿ�g3]���>��m>U��dJ��B����W.�I�D�b���L|�6eŞ}���`|iYj�(ͫ<֘�&����(�_���w��v���,	�Y�Q~��(!f� XW	xXW�Z�,�ϒ�W.{y��m-cU�JeiK����`�҄�����HZ!�����9�iWȻ�J�~%v%��j�R�ϡ���_��		�++q��34IX�����ȑWY��R���狤��^��}��Ϳ�s~����y��n�P���i`df����m�\"��N[ʣ:4��1ٔњ�Lsu���$H�:�HtqG����VK���!44 C��e(z��`DG�"ݿ�>�����T[�W�[��>�ՙ�2���w��r"��4�<������!��,<��w�5UU���a�B�LQ��V��d ހ������v0��u�[�#�W�߬S$آ5����Y���� ��q��@G�¹D�5�y�s�~� 8{wk�v/I��7��߾EI?�~S:6��.����싎��
����w���/�-��a}��"x���++Fȭ��h)�[�a�a̺� ��(�/����KGG�W���bp�M/x���]����tv~q�c労�K�D�jv�x�~���F�zy�������{C9�ڗU�z����5��q�@�|��Z Ǥ$A�3-�\��)�����ʩ2^
��l�xY۰�s�N�v	L����<��8�pp�JR�w/�Od����֏UNU��A�Z!!��������̪�qpX:�.>�;M�����ͮqŏ�4q�XY#��"R^�<m	��^Vh�J����������8_^nF�7::�'�o�D��O%�(��V>��}���7��<�z1TT,�{�e�81��COJ��uQӔ��\��r)�c.;���6�e�%���yJ���ތ��f�J���3폱�F�1��.�*�|��o�Xv��5&A�ץ���E�1BG?@�eí��</�/��Jk����}_�s,��^���8��3������W|K?���41a�}����Û�7���_#^pF��֚���KJBg�SS�3T��S��/��LM%��6������X�cp�������fNv;3�@I�bll��g�ڦ�����s'ڝ�MmD̵�<or�}}|� 6=��2;w�Ǿ��e'yee�V�^�W�5��&fiK(X3�v.�=��0���g�N�N����آ��D��z�WO 6���}�����=Z�́����?��CˤY] ���^s����j>��kQ-�1�֨l.*��c)�Qq�T
jRe��:�=���,�S�GZș%��~>�QL�d����a%L��l��<����!����ǿ7���_���p���R�:��:�HN�K���S�����?|�胵���Ԃ��X�?2�I�R:, ֲB1�o�&�ô�e� Ǎ�z��|���됟�|.qdTG������S��_Pp�.���@��AAm�Ifn��F"�ث7�C��	b]��m��gޢ��_.@v�+Gj�gH_Op`���u�.��J�출�VS�2}�8�L,�iM����v������2<�T	�iw)i^���Ʉ���W��j��)h�caaC3��f�::F�`�2sf�l��.�������t�u#�.��z�A�pz;z�C\>��	��z
��$�;�C�o�ٱ"�8a�7qV�	��$�R�����Ja���n��/��o\������ϐ�?V������^���q~qq�ī�A M�)���z;b����
�������ӯA����y�`0�t
c�SP����-OWw^[�3Qe��{`�"�J��$�ܒd�Fc�d}]��[���zp��\KK��mc�?8�1��@�43%�ڣ��ے�8�=��>uڻ�B��o�DX2i��'a?ށ�)d�HY`�F����/���N��L��)'���cC�I�^&��\��wojE`~�cuCU�1U�F_%$�#�~�}���T��s�
��_�����6f�/c����*��9�+�O��&��ʩ8ho����Y9{'c�F�{. ˩cĉ	�CG��f���U)`
��pt�zly����NN���e��_����l'3���g�zy�~��?��_t���9�	��|���²xEQ�ԤU�����9�5ܣ��TAU��d@^�z�x�d˗$hQ=jK׼N�b��c��e)!��܌Sl0�^4X�		��;���-��(�ww��bGب�p�޿OSp��7��յ�?|�����Zs���Aa�o������`za�M�*N6dyzC̝I) (Y��VMm��g�����k=6���W�UU�&���̆�a

���Uj#����I6��g����y~H��s�cTk&�B�fzj�Q+0))�����k�[��rsY�xC�&��?jU5�_��8	���'3�}�~��a]��+,��zu���PS�vS7�R0v�̯�~-M��!�6 !�>�W����4���ttvn�����z����c�T�~��}۫cje&"M{��X�#*�w2�����-�#y}A=���������ɉ�r΄�ݮ�>��4NM�~��탌�� ����s����ɢ`(w�,� G&�Г����*�8u�ذЧ泺5�%r�)��өi� '
��Carts:g��������:_q��m!@�r`' �I6P��+d��h��<��>}�+��������t����Y��7�E�5���11"%�����vq𮯵�7��RF����l(��j(S�tE�����_KS�QK���a"u��WW�[kVM[���C4�`ϷldB�=�(�Z��Ր�M���eږ�"�*uUU���wd�,(1�zZ����Wj�C?MR���1��'�B��\��=�bIU�Ṩ���΃��q�Im�ω�����Q'���2�[��2�p�?)�c ��?6`u���w��]��˚�H��v� ��;P���`�՗ş�E]:��2>�m�Ԫ�,��*�únp.=%{��K��P͂H>ū촠L-����	7�˗E���Q�znn��®+r�nb>o�J��nOV�tR���-�!(�s�+�"�˧AMթ6�_���{�&"؂�@�S��>���P$�푙�����z��H�
�̯�×n���I�J'�}��ͫ+�/Fx�^�
�n�S&l��n�7\��H��6�Hi���&|���:/�R@g㪫��/�����s��-�@ !F�����<�=��D�����P��k�H�f�^ֳ��R;Ƕ�?1���~-o(��;}_�
�T���>v��<��O2�n/�_X��������2���Yh�!�!�g�X�=~⨼���KK#=}���qs�ac���LS��_ɤ�m�:��.MX]ٍA����7+�	�Q�;N�^\��C�v����UQw	zttt�Q5M�K.e[�����r	x�{}��YN��<qV�������E�؊���n�ӡ��Օ,J��iP��-��V��*@���yy�D��+-�G\O�A�?~�(\<���:�SLL����ɦ��|*bL��w�.$8�^RS�1���B뾳+����N�����FsЉ���~�$��Տ��89݉��_���d%�F��w�������=���#��zt�{��VC�����Wf��[ڤ���V�xc(VO���u�����]��Ⱥ�+Rf!�g1�>I0l�hB��++�r�F�&���1Cm��5��A\Y���k_n���cyww^6v��O�������Vr��KS��9���cco\��~��w�'�uVT�TZX7��\����5�5�st�6{\JR)hE�����׳��,��w�� !/?4u��q9�|N5e����{����)N����/KL��~�=#�15L)�p=�b���#����_���1���w�\�Y�߇}}��C��W��]Op�����C
D<��:�2�����X�8x>�v�UIp�8K��/*֫�R�y鑻��Ɩj���|��ьs�3����8޷8��������Ƶ�ͷM	a��(;��ыڣ�C�α~�춴�;��B�2tW�E(�[BQ�T|ԥ dd�/��v�Xֶtju�9ܻ����/X�uy��Pw�D�-V7j] j�7t5��1����J�]{LqTh��9nh��{@���#ǋE==�N-9��T�=���o�W,��Ҽ��Z}Q�@N�o�ԃ�g'3�z�S�z��� �m���7?��]A��-��5dU���gD�J��Y���*�bw�'�
�G,��n97t��[]_]�h�x�����h�H$�fu�.�Y�n�@EAA���}���?���4_�ژ���o��Qbv�z�ʨ�2��FˮE
�����_����ffp9�-�m��|��07��SL��������AO��9>�8"ib����u
\H_O�d�O����g��7gq5�L0n*V�"�A'ʓ�c�O�'�펷{�]\�����b�"�XG ��6�
#�(JT�oK�ۏ������Ur�[�ȫ��%�i�z���B=����J���TI�d��ex���ʣ�0��7 �g�rOCuf$%�ç��dT;�g�SO�!��^X �G�/�L ^���ۑw270`�\���ս��W�Wr$o4I�������V�V��LISe-�adU����Q��POo���s���y��B}�S5kjy����Λ�7����ш`�ϻ�ω�	͆���/���Kc-��CG��OǮ���2 ���u�yଇ��P<��c�â��a@��F�SBA:�.��{�n	i陡KRJJ@J`H�i���3~���z�d8sf�}�^��Y��x$3��ƅ�v�W��R�ߝm3{��)�&D��k�RˠN����[�VK$F�'&�|LL�i�?��d�"�E�w\Pk�z��]��8�D{^!�g��޻����K&�?~��q�a&ty�S�Rh�f�y �{�ط���"@�vx㯚�3�hߐ�-.�cj��ە<��dh ���7XGW�AQwX����r}Ԯd^6�X� Y$���c%���>&�J�7Y1c��c_y�p������K+/��rc#������r�/_��6��Dץ�ϼ<�i%`A��	T�^�|������SK�-a33����1F��Ce�5Co�c�A6[R�t���J�8KJ"Z�� ��]>�t@DS�l��O�/_�{��''�N�Ճi
݃0�1��=}���n/�^���ί��	 y�$5]��z�o�C.\vsڒ��Ir &lho����WN��Tz���DP:;��Բ�HL��}GW|i��{��a;y�1���5�@f�)��/�˙�Dy}Y��'���Y'{O0��T�1����Q^�J���v�잭��.7�V�O;3E�Ғ��SRE$����?	�8||����oɈBů��fy+,� ͑l��؝�%�E
1�|�of �@�������BiL��T�ZE��3��C��g�H��5�,���mw�t� �/�Wqw`vtt`�����~�����]����:ȅ!׽3��� ���qk2�'Bִ�bu�DG x!n� �P�H��W�mmεX> >���v���GV�	���(�imSq�3Y$F�S0Hf���¹8ȍ>��װ�_����+�`�LR�����rqj�S��u�߮n�?��K��&������{]��^l� <�X�i���f� ��0�BkV�I�m� 5j�����k��f���)�d�JŰs��4�ZI��Mc�w9M�|6��O��ɉ%���t�1��J8��B�����Ճ�4�̒�z� �Rz+x�*������M��-8��Ä݃_���Qȓ~zw6p�'���N����r���x��I�^������TC�8ş���o�SmY�T�Ip��Es2t�5ǵ{k�V�v� ��-���;���pg9*������L����^P'���=#/Fnott0��]��m���2�q�f������]�5��8	�9m#���b8�_�Q�b�BQK���+�~.�u)� Fٽ�bs����uq[�֖������]y��陙������d�J�'#���a#EA0���Yt&��*�2 �y���b3g �{�4��X^Q�����2ޒ�GR� � z"�V�fDଘ��2��Ys���eL��1�x50�[�-�3z¹����f�cz�1I��?r̩C��c�<���r� Mmޑ��EP_3�$�y}Ν�����H�n�)�,-1YR�$[��%��*��(�ק^R�!�^���O�	��v���g@���y�/-��{/�����!{%����v[Up Fݝ�h�_����&Օ����E�oǮ�ΞN��������G{�� ã�	-׊�c��(
2�?��5|�����K�,��`�����RJ��`C�s$��<ʩ�J7�#)�o���;��Gm
/��2(̾�~v�86,�2�E[�nň�Z���N��+������a����X�K�0��eo\@�>F�Pn!ߗ�+Z�\\��'�0��{���Ī�c���~U��B��(a������N2Ʉ�^�{Ki�r::swK�Ϥ� �����.M�\��oݣ�_zjk/�3�o$tu��Z5O��F���|3�+?o�1z�SPYI��l�&��j:���LM=T�
���F�Z.ݔ�b��o�w�6�2�'�����M��#,z7}�JKN���y�*�M�n� ��_RT�OY�+-uչf6��"H�hG�a�x�g��0�URTT�"����l����n�������t"�v
" (�kGK�҆d����Qq���Q.��.�T=7��O m�!���v�u�9�c`-���?�LG'B����ܠ?"\=��C����{�h��R�,]��e��	/X�83#��)��K��Y��˾HN,��_��`�9}�SQG(F�,HC���,��*\��#]��Ƒ�ƛ�~����Z����-I���e7qb�W��,�����eN�,F:��,��˧��Z#͂����R�<N��\�aF�󹧍�J��9�]I�BZ�1>W�ꯏFR��� �MA�eǊ;��^|�̋/�ʄb?4���v�-<{�Ì�+�������܅�P�4/�~IC�Y1��KA'�
����-��c�ΰ	�H.B��`� pÄg��)=��Ë�St�E������f�c�M�#�d���l��e��q���b��{�zt Yl㓍�W��2W[LdN���Y��E�c��N�ܽ�a1�󌇗w]�M���MUO	(?�2���6* �SQ���MI�JIh�ٯ>8D���D�{%�>2,*�m�9V�m�����`(����i��l*�����������(1�Hl5՟���lr�mաq|��w?��}�,E���ƋY=Ҋmm~G 4P��V����u�����Yʨ��Gs_-�U����
��ாã��%A������:X��0]���DG�Ն�_�%�_	@����n�:��4��A�f�E��ID�w����V���T�[�F��9	+%�eoBj�!
�+� P�X�_
�)07 h2M<y�|Lf�"���7p���R;�/[��\�l�r|o��.a�9[Ygn����f��et�����|N�[��t�㓀�ã�ifF�9�Z���5�֠x�	aػZ�
	$�de��d�s��O���I�fB���j�|��\�6���1����N�K��$�L(�O����y������[���X�2{��E�*�W�%2J'C��p��Fߥp���3�j�q�囋G�{���s_m��Ct�Qf~��"f^���K��A�z���+͛���D���l܇I�	�jA����ǝ�?����ޘ`��v����@��7�Ȥ@�n�������y��}
?DC}��RØ埀��9����0�����mE��F*M��O�^44�´'#"c�k��E���I?~��쵶J~��`���},V��"}�x�o^�����V{��]�X��)�/q���O2yN]0�n�vӸ���WΆh��eSC�2jh�`���^���c��<X�8�2���wȟ\s���G�K��IɠF�+ S��E�__��5��3G](�9*d�3�Z� ̣�%�8������|����}������=�с�(!�O���K�cg������ԥH{Nw��eP���u^��'C��M _��.�65e�������ֻ�u�������T%��ܤ�� ��/+��{�߷Xȃ%{��_ ��u��ڟ��m�{�:���ʽ�����\�#:�=�Pg�K�1BP��`�k����>�6�ujmK�\�����o>��%�O�Ir�Za����d����n��ER���ÿ�2���{S�ኲ�z����Y���}U����xj�5�Տ�q3�b�~���+64>��̤T"�e����wڤ���$�O'A����� �<�p q����a�6Q���EP���r�x���4�F�yG�8����9H���oN�V��f���%;���v�/�:>222J�͌q����y��M	u����3�Ya������rxt�X��Ž��D<���1��4ZX�Sy���$��&|J��1v7Yf:Z%uׇx� /X^^��b���F���#���'��#ے~Gg�`u���'�8��?���*��QZ�O~� �������m��w *U*e����m'n�g]���%��u��2O/t���7���$$�	B��_�F�¢2oR4�a��ն�����S�~~��w�~Ql���O?�
��䴴�LƤ��G�1'
X�ü�E+������' q�d���1 ��U6�f�1��;1B�Z���M��»1�oz��6���%���eâK�w�üJ��=��*ݸ��N>��|�������^��/��$ɜ��!��%��ZD$�] ������Gz�$)��j�����=9V"yJD	y����g]�!�r/�+&���L����	W����XZ�v�+$��[��1�˞�P���8_'׊��N�^���-�6H��x����a-��0���k(5*}}����ޭ��<9�$��Ņ%���zc���|b�m���Nݨ�?`r{�.��K���~����k��Z҇�y�w%�����_-.M�����rw_O��&l|]�3xճ������ߣ_��I��<��]XV���e�]nGG���e���lM9{���|����}�B�4��_��o.���H`����9^
}�_߳V�'��ӝ�'Q����@��кz�NL�-�|���=6���8<�B���-�[=Q��4�y�2����[r����΢��P�)�^6�Ք��E�Q�("09���*����&�"�x��	&��:+�Ϲ=(�+�h%��D�+���|O��C̷^�QJ��Q�>G�2M��eDd��]Qc�5Ӟ���B�\�� ��af�n�
ӻ�k��v�aJ��o���4����*�����ڶ�:�,�~W�%3,�j=�z���?hoS����
�cd�SU��+u���{�Q�7�Y��pں�������n��<�>��ٛ��M=�u�4�4,U�z1vZ�o{^d��1�l|r�V�6!1 �l��<='/B���j�+�����3��d	@$1I�
QP����?�ݣ��H��;0�̥�)u�9x�=��z��3,���kC��. �ʆvW����"�)]ט6`!]�� 	Q�|��I�K��K�66ۙ����<Bq���e�>:9�L�M|i�.b��`����wsE�o�{�=�89��3KFZ�����@��a/�<DP��.���n�(��J麔B���9�?Do�~��_h��&w";Lu�o.  ��}�+��bt���LOd�	�p��Tע�۟�Utx�r?$!�rq=<̂Az�Cn��:����wwH~R�bع��i=_#�1$lx�@�3H��$���q��� ���<Xm&E���O����_i;.��'og��A��ݚ=�+�vӿ��?I��e
�K��|�j��*���J�&�9fj=l4à���;k++����zt�=T	]�`��D�X��T�N��Ǹyw����HpC�\�Fg�9�!C_%�le,&#K��^rO�{s]ή9��q=16i�oҼ��Vk��NL�?�Ԍ��g�����B���_�4%&F��][��n�fD�%���xEE��D|8e7g�Ҫ y� �V�:d�gխ�;��?��E^�.�E�����5�U6�|���T.(��+e��ڒ����:^~��\-��=�ͫ�xa�]fF&�WGqxO���[�Q�����x��b;4��u_?ӹ5�^�y�Sʅ�'�^�n\?�Dk@wH?~�mfY �fi��e����uO]���T�>b���������C~Y3޳g{"�Vc� @���֙ys�V�P�ϽQM����ٳ�<�%�W���j)8�
	l0 &�����Pn}t��}GT���V+���Q�Z,���ǩ�g��7��ڎ;_�/K߈����q�͋������<��\+y����[�L�\��D��r�ܳ�M��:#��!$�/<ߕ�_X��yc �O52m�ύDg��.�ߎ��r��-,J'�.�u]4��q�|+�TJQ�6�ӧ��_�JJ8��¡���Q^hԇ2�?!*	s���v���d���p�5 ������R��T9''�I�ȝ�iA;;���lF�`|\,��g6�H/B�!3�<k���,=����r�fi��F���%�)@����G���1N���Y��JĠa�U�������
u�4��d�K�w��uR�}M-"���N��g��,���C،����X�F-���!7NYZ�¯_���}���E�N;�[A9�Ԉ���V�^�+w_s#�ȉ,��>�'���\a`77X���i�>�����G:�y����ѷmo%a�l�AX8z���.m�������F�Jⱼ]���7�3��ü;L貊���@�:����,�0	FCC�G�Ԋ[�ȤJE�'BA��N�v��6E�Dk�F��O �Ԕ!�'H����-�m7�2n6;�
���F?����nY4����d��#R¢s3�	�
8QR���v���ҧ�ߓ�Nn�uu�y"�}W��<�$=�ѣ��IC�/�x�'3N>8F!G���;ĸdI���R�&�2��VI�Y�W�^�m���r�73砻`I�WZ�����s�%-o�Цܨ��!�c P���U@���~��z �"�E��ϟ��Η���F!!�W,Ph����$R�_���륙w�Ϋ�ڂ_r�9i�!e�8[PƟ�D(w����H��=�rU#��w�;�Ɲ��dڄ��*5�;��(��
"f��nx!*AqM|$�v�I�����M�Y��.�;�I9�L�,��
?G�R��Gr����R��UTW��«�2�f6�K�J�"̄�5_�~�H�r�k|��u�g��շ�Ǻ7�C]r���m�g��9�۔��]�����`��Z�%a�ܓ�a �1I��@eI/ԙ�q�P�OEmm���t�B��4�s�Q�V.�����$萮����a�*�� .��M�$�zIK�NW�̡��l��< �/qqqsVժ�o]�'q���luaQ����� {�����J�9�|=ޔ�Ae}}��g��QieV�7�~9��w>��r��5������1�j���?�O�I����=�#iv�g�*>s?�:9�S��"��1�K��$���>���官�����U\<i�7����Vy�E�C�bX��Ք�<[04����j����Ȳ�HK_;v#],0�7r�1��ڤ���hT�WL��H��w3]�&�s@kE����4�^
��uq�g���� |�mq���s�������/��$�m���Ft�2�6���\@�����5�A�a�jMUy�FŘ��$-N���ȅ�->/e8��XZ��?�;*B�W*�.|��g>��8, fa��8�R5�?���F�[����F6=.��a���lLr]��C�	���H��fG:Nc+7a]_��7�$-&�������VvO_�Gh�u�]8?�E����M���OQv��U�lף����*�3!����\8����C�b9�&wh�ji��$�	��������Tnk\LI��'(����o�>ڹ�Q�xXZh��9�*r���sI֫�qj|-H���Cٳ�æh���Z��X!4�i���?�H0y���:2�ի������5��,X�lR�����"v�����2̓@�in5����ѫ�䟌�
]a���I >���$y����b�6O�"��-S݄L�:ݸ��5�/�вO	�~�[���(��H;��d�X��(�m��%q��u���+'���7��:�TP��u��#$���!�D����]�O�����<܎���p��F�*��E�?��[&��I^��∄���%z�,������Î�M�1RU�}y(8S!�!��.��X:xAl��1��1�&6�c����گ�|'~_��
����b��%�S���)��=�O.$���\y�F.k�\s��~I�������������LPcCs�>��![�*�b�s�}�B�h�D95�{�_R#��
&�!aT�\�nu�;�|��su�))�D_���r&޲y)]^���3��.������Xo�
|W8-��P>)h��ͳ��v�>�m�j4�pd�BA�ؐ���d�:����'�S9kEsƆ6]��]�g��R���d��6�]�rӵc�>,,�Z..H�+u�	m���֛U�SU5�>�zi�1��%���Jܦj��x1��s}ܕ�v������r�ۮ٣��Y˧���XX����y��C3��;�mC3�1H��c!�K�RP���3>:z���7�66��{�j���F�ҳ`��(B�ԟzNp�x�O6�d'Yq��k�x����d�5�!�𘿿 ��Z�@��t����1��M����)WcY[o�������;�	�*��6|�	�0u����$�8%���;,��i�ʹ���߳�Q����ݸU_�N������z>o������\VZ��2�zK��rL��m��Eጌ�7�ܵ�223Srs�&�1��J%:�%4����Ǟ�Lf��ξ��/0�˹���`[�}����I�C��dvnn��M�4�o�h̞��ǰ1���yu���~U1��"q�*�==��8���u��0�f:7U&�4��y1�B���/�NF����t+�U�K��}wجy�i�Nee�K�ehn��˒3q��[��Q܎N�C(c*�Dn�\���^WL��	m�J��6�^�e���a�0����sXƏ,?qm.q_�y­�O�K�����7_?��L�<}�y͌c��s�.�+'�;4
�#oY����`��(�׃�ttذ���������h��`��5�M���/<��AjS:����e��wD_����y�e�J�v��e�*���
����n݀C��CKu���8pqo��<>�M�V�4,f)�T����Gn.N=��?�KtDr����j~��	>��������k_�͛��7?��̠�H�B�ԩ��O�g9���0���d
�"D6�4�W�"S}|+��A���(�-��e��T.a_�K�W�H�h�����}���k�J��/���3/�f��3�[p�߇1��oc��<<���+��kb#8�r_��*wK�D�ٳ(�XC>��ቩE��^D`�j�tFF}��766��r{>"�}�'��}4��n�@O�9,�s�y��+��i@�;xja�U�i����pfF:(`27��ߟ�Ye�Ζ�(6� (l���I-�1�����$p''���/�mq~�� �<4���h�nN�w�-.;��U�Cimb^�zE�1A��ͥ�,�S�����f?y!�y�M@{�ų��AQeU���%���j=����u|;�#H��D{��%2����;.r=����:��9�^����R���<�<O�7�7M=���I�f�:���E"��z��Rpn����92t��9�⩵���������}�����=����c�4�Ǔg�q�e�P����2��=mmm���U���E��� 4v�4I�.��&2����+w�Fg�&���sG����W��g��NNj�9M�@���?!|����Oz?��/�|ڛ􉑫�e0����nd�ts��%:����k�i���r&"l����k��d�Ň>��&�V��$MV�yӌA���_���3���=�g��b,Ȼ����q�ߝ�Xm�]'�HOC[c���[7M�� ���/�zh�z������2���ޘ'Vtd_�|Y(���d�^�,R�����q��)]:*ҽy%��X�A9��{��{z� ��L�.\\�S��{!]��G]y��/I�Xh�§�Y�K&�gRR���'����kS$�e��\t�ep�g�3�j���dN��1}�y����G�D5�
Ȍ�ݨ��M�4�cû1?G<���"��ty�}��O�ߒۧ�2�z��H�=����M�J/R����q�s������#����P�`[����[t�ϲ�l�꭫�ka�7+d�x�.����7���m�����bihVv���5�Y���R��Խc]JER�O�M�w��I���	7)�^(N��� }�q���=�P�0��؏Q��י��,!�//��RA���j�tY�X���O��y�aQ�������1�������$�]�%�Gվ��u{�/i>��2>�<
5�N5�]Ye���{�����W��.�	ܥ�}���8=�]���¢K�������o"c"�24Tظ!���8�D/z{G�e������G�ʪ��^ǣ3XzN})Y�l��7��}��\�-ѭD3<��f�u�@�I�N�p�e��^TTԛ��|D�ldԌ�B�QIt����Tr��o���G�����U�Z�?����v}���jeNӵ��j�u�g2	� !�U�sݔYm��A5_�=sä���^�Xs%���XX��?��?��e����Y�P�LP�0������)M��Ov˭s�|,  /�|��z�w�,���w'@��:X~�0?���]�G�u���(G�����hK��"�+��]���x��0�n  �c��D���~*VKQG�,�I�6��ۻaL�gA �wFu<B��5a6���2{?���P��� �~7��[�|�����ҾGh/�����;���J- !/�z��f6���B�P�a�c�<��i�Ǻ�J��G�����EEiW�y��U��=���CU����M)*t���bN��a[�ם���C����z�F�Xރa�|�8͍l�L()3-�ߊ�.hlR�䳈����]�A1t������ ^���E�'��I��^�^p366����yͅ>��������%�H�)�9��e4:
0���hhm��ee�{���̌Ho(I�jH ��e ¬���ûCSN��T�%��S���h��+��MfƁ+��1��'�qg���Y7̏/��A��>"�p ;�]]KK�Y"�rC�rS}}*!����JM�C�LI������$3����k��<U�f 9�<g�3��ԫ5~��䍒�毝��MGG�c.��<��WZ��V��gkPn��7=��B�	�#��M�". ��-.8¼�v��֟I�Fq���������[^1��/X��� D��	\�����������⁅x�*6w(v~Y*��b�v��b��ckW�;�l�������Ltj������O��Ҿ���6nS�t�9��k�����m>|���G_���0p��������]�cK	��T��-l�����}}��>�?�4�k�wG@`tpqRr�$=�ÿi�{�Է�	���1w�9����HK����{��#b�F�j{��mݢ�K���߽+,J�_��s,��O��DM���#���lo��>���4!��㾟��so��?4c�2��JAȞ����`yٴ=���n;�y�u΅@��N8(9j������>Xz��J���!�5���A�`�[�<�+�3����ˍ�R����+���/μ����m(��LM���8"���{���Rl�Z��j^�q�ۢ��B��}DR�������4��9�Qk���Y��^0�H@@��:H��҅���P@B��*<��P������y�HEUs3#Ee[NJ��Q#B��ݵÑZ��9�C��d�:6:�wv�T������ Ox"%E�a���C7�*F�w�b*L��������m�b{K1�1W�vĹ�}rQ���Y\&"$�h��s=l�봖�	�ڴ�\v�S�"o��߯?]	w�_�����o��~�h�>Ҕ��~�*���Mη���o��x�Pt"!فYŋU�5&vkK�kc�Q�T�����йAUC��, R�Ҽ�6���-���'�DPS��A��V�0tZ8(Y!�W��3v~��;�޹i�#��;��Ҳ�Z�,�Åb͆��G�3��NB��t��7kW�d	*ʮ��k���'嗔ਥ�gH~]�\g����zd�U��MY�\괁�x��s����偖�\,{���Ծ��Dۆ�ab0#Z�I9�yބ{��F����C���,��H����["nHe"�JV����7�������g�j˒���5k�����H����I�~��� ��������ggJ�z��$x$�%�=���D��l����$�orHM
u?p�0h����ǐaBt/+�h��#�H�˴-Uj��R��=Ӌ"l�pC��\gr>�;���"Nr�~H2���Θ4�Y�఻;�����:&��> �n7#���<�����s���"���;�?�oC�	$m�H�_W
�%WO9i���ӭ��{�䣮�`{���?!�3?cs8��-`�U��(�~;�Go�v7b���Os�T�����11�UB� �a#{, h��bR?�da��#'�8j�v�_�cӥO���ǏY����/������,H#�DZMbj�3�����(�r���&��\��H̽��ѓpU�g��}Xe�G��>��K��k��j�~uzIO'b7S� D}Q6QX���=G��U�
yd@D�~0遀z{SQ��)]�*���,N�2̠KeG,��5e���H�yw�{'��k��?�z7"�X����J�@��Ǽ�!)ѯ��b�%�9�O�.Wg�Ǫ��p����!�R�y��{|/�~�Zk$	�1�ϩor� ��Jک�K���ޜ�ަT�+֡�ܒ�/�3O"5��'��]mmq�,�^�,M����'�l,c�.�K�#�N��� `.�6O�z�.���RRjQ`r;���;J"ʏ!]�:%*����!�H�(2_����.%e��Wp�ct��Ό<�3�/zf���#�w��o���S�=���`��Ə���D��q1O��d)��(�@���1d`�s��p�ј>�����1�.y�A)�i���pH���\���L�}��%�D�����HeyD�%�,����Β�tJ�
p��Ƌ�	־c-�W�T�OM�W�ƕr��P��~�Mljj*��TP����^��XYS317ri[�=�W,P�5*щ�>r�����-lh�sw4t�(�|�F�6��4#�t�C��}�	�J�8���7�h̕��[� H���6&��]&��m�4����]x�<1�)�P��)��٫=ٽ�~��+R-YdIII!x~�A����щ
a���l�� s��6�!r�c즐�&��뉼xle`��*C� �W�u_*��ěEoaq��R��@t�=\XXx4v�ĀV�n�u��t1�88|_h>Y[�kXoZt�p�(E�.�H4�y������L3���$��[�˻bDp���Y�lx���qP2��	6�1��@H�Y��Q��� ��(��u�-y�2��	������l�����Bųc1Q�r���PQy9��'*��%`�*�/
�#a�� @�uwc�Z2���ȓJG7w5�Y�7�X�}x��I��,�/�VBk�<�w�Ac�AwCܿ7zp� �_�ɘ���\���c��u*��%ps���ϕ�4��mG�>S65���|��x��%���Nll�Z���14�ot�����Il�+*J{c#���c���ܿZ�V� *%9h�mg0=�'��2B���}��'�?ub���
6ŷb��C�2j�������Fc�����B���/��g����C/v~i"���#�ן��}`&u���c:�)Ĺqx�����R_��U��| �;BD�7$��<
<���||�<�P���"A��������]��ר�%UC�B@H���?����՗�����i��a3�;������:#e2H��eS��P��,���/�N!�����6|��'��(�@�b| �����f!y�PS(:8�s{�[�Ě��v�����"ڠr�j /&�E�\�icllllߐ���!Z��DD�xx���� nj�I��֌.�z��H��	NW��ר@��&ߐ��W��nj�?ݤ���w�F�q��s��.��͑7_�ʊ��Á�充8��|{�}���BB��r������ܜ�ق�սW�d�}� �c��h����	�x$,8qV@!�f|a��wP�Q�Ě��1��4%��H�v8^9�����V��Т�qll���@�84G�1����a�e����-	���d�yY-����T���:L�8�z�sBqP��b�n�4���7~+�����[��'5נ bW8������d��Ӏ&SL���/M�z�@T�h(k+/9�8���i����ə���xUa,�\���{o��b���Y��������S���eӗ�gDD~�)�)G������zN��f%|s�����Kd�����w>W3Lů��G�EE���*���X����Z�N鉉�?,,��"�ۓA�j���ϓ�;��U�2���WS��ZY���E�Nx�5�4Y����2���ڱ>���D�2����+��?Ru�[�Ktnwr݅k㸡߮75O��C}���\�ܪ#�Ɗ�#U����p��B��$S���"`��E[ftm��I�IS�G	��چ�x�j��
�\�ɒ� 77�����V�dA$�&�(��� +OfBԘ3�"�[+�f�A��վ��O>W~�pu�OQ�E�N���z8�����ގ�a�c��^���.��/ �Vc�E8�C� 64��Ck��K�j�4�ֆ�<ڗJ���v���E2�D�#w6�3p�mٞk�'�~x�8dwé�Q��" �$���M��N�<�t�z�㦭�_۽����-�?rZ��_��Wd�`^	y�{<&! x�&��*�#WMH_joϑ!�/5����jY��zo���d�驧�h�^[ � .N�O��������'�\���٘�%�(0�LK����w����@�&���~����/K �}��8���2f���ËC��HI*w��,'./Ta��lfl�"
�o(h}u���8�
���0��APLP�8�r����+F� �q����y�ĠZSQ]�s��߰��J�A�gq�KƬ�X����0�S�7�(�EHFy ϹtB�KS�"\��v���ҌW��ٵo^S�EKSx�f� 	��KP빮�v�S� X�9^� j �S	Ű����(g���j��~9M�~q��h��uQX���瑹+�)��c���:�).�-&9o�M����+U�UX:
�#�����'��ˇ>��K�V�M��o4���{gi�~�C��L\ۊ�pps���?(EA�I�?9�#:-^[ˏ�,��鿠�C/2��ߛ���Ʌ��%M�����՘W�f�������_�^����]���P�F�%)H�����w������R�8� c���ws#�T�����'��w���l��|,b6^(���le�L;�B*[�ք�wwC��y�z���P��z㛔:�9���&?��j��r�l�
V�L���`z�Q����q�o##�3�o��$�o�}���WU(�O&D�T�b�?"�4lj[<�A��ӓ��{ƫ������7�-�j����_�5 v��pZ
\�`�`fz���$�������o�x;>>�R�����N�L���1S|�������8�/����,����nO/A���n�����&+���tM�ގu�`#��% ���3���j��^�>��!�$NK���9���h݁���Z��덦Ft��ߗ�1�L���'?�k��y�k�d)�8w4��U��T"w/m3�M��C*��T1rkk��b�-{{��<��F�O9y�F����htt�}�\"/ˢ�yَF!�ݻg�S;�4_&����~�	�N_��џ��0p�,���)���y^)q�@�fS[���b���y�OB1�n�"��sa9*��c* a*H���5w��m
���9�o HB<!��w���0�����"���*�6@I}Vz]~�l�ˌjj����bO	����. iM>�Kؓe#v����K(]�'�S>p@���H7` B��%�\Y���ػU�n[}/
�s�F�m$>T��q(�E��]�����M��:�/!�o�W�?|��/����I9}t�����C��46�P���Z��P@A(���x�5b:;�@�$Q��-� �d�d�&�O����Q00�*0�7fF�{1��%$����<�|n���BL�|����d#)\r�H}�̴���\lv-q�,SR�]C� &s�!?p�P��o�Ȕ̞���9�����s��&���o:vz$��¹��
����$GӀ��\�ѻ/M>�h+�����y��јd��.h��e��M�CP�b��#?�ϟ?�?�`���1ma�j��#E$�5
v�Q�Ve��--;����S�F���t��\鄃^q�f��U �U6E��S݇n�U0ɸ�I��N�Ǫǒ ��c.L���͙�8&�r�o`�?��v̷�������ivc|�ٗ�V,F"������UB��h�H��������B��|t��9QeP��4���� U����I5K�p�����EOdݘr�C�ȝ�Ɇ�z-m��w�+�3`A�=�F:��6���IM�il`Z��Â�|ߴ����`�}�9i������������F:����bs�ͣ��RB�8(����N���NyR�/G�����u� �횻7O�Y��:�f@7�"�ry�א�D��?�0g��K�}I��B�EEᨲ��W?n���V���˦.�d�ϝ�Ґ�Jĝ4�e6��ɛ��VR�bGL>sz6fJP�I3�V��;<<��`�1ou�t]�kQj���ݓ�I�E�����t���	���jnӲ)V2�����_��k�C*��k�9Wo_�^��)Y$����h�������f��h���xCj��>Y|_H�ڨU��ڢ�J��k��%�r��������t��\��%n�� q�g4Q�)� ������
� �򚚤;ȝ�o���^��ࣥ�iL�8S�� �4������*�<Al)���>GT�ǿ~E�:�4�0a�[�)+p��1��C`��͏�#��
�b�Ȓ�\����n��8�p���i�:���ul�oy�*�K�
�󿐠Tt|�
�̀��[1�.OSQ��b�+a��%� ��.��	=���o�����]A��5?6,.�V~�/�?��2,���F@B�������QJ�Ni�))))�N����a(�!�K��3����ŧ��9玽�Z��B�2��\�����5�7��۔.}5�4����j�(�\���i���Fu��[�ˮ;3Cܝ�f�P%S�Ňc.����1�n��N��k3P���A�L�)��~6,rǢ���t}����Q�&���jT�C���=C��rn�����u3�Y�(����t�}}}r�sXh�
�O||�Y�"j�8�=��q3�J�r��qD�	��|ޭ�7.�R0��X:`���vsä�k��C@ի�oC��N0f�Z���Q~�D$�Ӥ���]4W�Sf��ס��QQQ�����/��c�Т�_Ih�_|\ڊ|΂=B��J����A�RJn��Mθ� �X�rS������7!�s���`b�KQ__O���񪹸B%���}ec؎x5�+�&H� �M��x����c�:r}w��M"��������>"/8�,�3$�+�������s��h�L޺�������.K����7ֹ*L���	V�(((���"���r/]�`��������c۬�j���M��_^��K��acc��u��[�&�c�D�'��Ե�8�X��k{��d��AUN�����N�g���#Bv|��l[�%�j����)�ʃ�^�[�����}�v�xӼS6��Ҭ~/��g�+��$�g�n*��h́�i���A��2A���:l;�G�!�# ��=���0*�`7�{�l��b)f���J�8jn#�?��h�yd�Fs�S�s{�C�����6~��=Qၑ���n��@
%�
�9E�S��||>�򜁩����l�	
x��*(��8H!�=b�S���D�~08�1v��R$f��U���{ Sj�;�9]5,���d�%^͆lnkp�|ʞ�vOC��]{���34ć$QSsb�mVVV
��#�Q���� 	Z;{��y��s�^%��t46�?.&�� heq�n/W��>C�m�o�ɖKV �T��~�ׇ������ F�$H��SXe���IH�j�1���V�����7�H3H'�y�^��(��tjő[�477{��Sb�j�={���}�u3?d�E���l��詙�q�_t�X�j����S��/�92����W,��"yp��(�@��o2��qn�q&]��go��:�eao�mb�P�����碎g��8	WOH`��T (���i^s�R������{s�Cx�Q7�{4�)���:d��eˬO�d�g_���!�X�0���p��?��7&:��	U#�		��)1R��w�=�_�g��?;�7s;���`���HNN�+k:t�rq���QS�,�Vg����5@��,*��l1ۼ
2�k.�. ��؝�vzv*p�
)��I��y:"h)>��σ�ݶ-=����C
��+���4���!c�c��#/?�d�����
lw��h���*��t�۟��C�_�D��J#�m����ϞA HJ�H>	%kko�WNp5�PS�Y�ARۅﶌ��l�	%�q�����P��cZ���{kI B��� ��o�7�ʎA��֥ʲ��m�A�.�
�?q2��mPhRRғ��1��
��3��C�m�zSk6���j�_� �փ���?mϘ��Pm���0[�e���+-SR7������o54������Y��,��.��+x����K��q�9��������"Dމ̒��.�3;^!��e��os~�>'�-�o��Z�v�����3����mfƖ���h��H�����87̓B�~�	�8���e�t���kB|}�����-n�0�E�����2j<VNVY[AJ����b��o�E�ӳ3�
ξ~�b����g��tv6��u2��X[�H bF�)�[��K�#����Ҧhd@Hv����7���q����מ`��mQ�v/��X�����GEMe�\�L��(�GE����-ZJQ�w�5�u�����`C0TJn.��j�M>�.(8���t�W������
9Hd�1׽��FV���5�n��զl㞡���6J`=dQ�!�X� s&�A���Z�Oqun7�\d���J��|���6ʻ���ج�
ˉ?�on�d�W��������Qۿ����g�C H�����?��5�UY�3V�1 �GG�ˣ!�����+��^��ⶸ��=�ߋ$%�F�(�w����4gv���p�86�xw~�#0�Y��pr*@��P�/��O��W���<#� ��ӏi��f3���f`�哥�;����ՙgFG��D��O�,0�0ao؛�	^;�gS;��#�Q�:��O���#�k#�� �"q��ŋ�T��Яc��az��C�����'I=�X� 9R�[ �I]�r3,E}���K6f�sK���++����O���'��T���IMK&�kj/J� �<�o)1�no��D~OiO.���H��pqͷ]���I}2�o욨�щܙx��ֲ�AT�ܥSr�곳�z3NW++ڶ�vE� ��W]�m1���Z�+2`�?8$}���Q�mB�UX�l�c�������������LV�y�z/xh��̃�(�[N;PLD�l����])���8}���"/�����~�����W���T���|--�:p�q���"�ȑb����^R�1������D<�'O�n�B-n����g��l�q���2�<�� �6���o�¢�d�^"�y�6��z�����vd@��y�����, 9��R���QH;H��' �
���9��.s؎����oh��̝Ԕa~{��R�_?����b|�|8|��͊��+�]�U$s���#��>hw��zJ}��A�VWO}s�UWW/�t�"|�T�����
������S�z�8��# ���4�z��P���Mg�؄�#�c�1����uS�������(��N?3{�iݳ�c�Q�]� T*�����EF����΅��Ja~�`#T"7��ƕY��Mw:�����6/99��\m���س��en��'�:#H�EׇΛ�_�)�,!΁����g]��jI_�I'FFƉ}��*��I�fO�\D� v��P{)�$Y«��W"݁[�������m�"k�kH������%��R��9o��C�W %NI��4��z�~������t_�7#I��"�I�)N�B �����.���jmiZ�1`o�6���vu�f+1I��/��}�\GC�����	��d�ކ���C�wHY��ȪhL��ҷ�������=殀������
�.d@�wOYXzW��p�[z�M�A�+	��[ԃ�¾{3�NB��'���LOq>$&ِB���)��Ж{�qKڪp�b)V�l'�l�k�oK��fM��/��q;�;,E�3�����^��!N.��~lT�'R	�A�n_#5�`e��S��"^11qP+=m�m�Hp��br��u7��DIU�����b�j��t
��s�7<��By#����T'��*%�N��qg���l�SF��p_��gs��?��Z���#cՑ�����s����X� X��q9�⛣�Ya3
U~�����#���^��x��/6.�BD��
�U�E�����GA0u5`?��~���jz��`�� ����X�غ����J���V�r&&'���9�'��r�(}�,*�S�J7���I�>t��p��~̴!�դ�{}tm��4��a���������s��z��ar�Ķ�gb7�$�5�ٻ𲟱_�J�����W����ߢ�D&B��vuAa�2%����I+]V�3�'Vꋋ,,, @�~�ͽ󠥉�%��UН���c���sL��?"�8�'��Η�)Jj�!~����\�Ƕ��|kk���C^1 �6�\��١�����g���:4꼖��v���|t��"����26��BUEX�/�q���`�pߥ�b�1�J� ������;�!!�k���x7GG�ƨ���?���3��_r�֔.'Ҫ�a�߿�?k��B�݅�"P4J��`���M--�)߿��*�� %�����UT�DYU�?�&[5���z��D��<��m����m�"��@%�d���w �jmS�:ۼ��ٓ�x��?����E�+Ϗm	H�ּ]��SzzTm-�?�]�,ΑI��k �pi���~��Qg��Z��$�((^g�v�R�Y�7_��(�qL��x/�����l ���S�E{��FF��g��7�垦��ڊ�����;4ӫ[�J�vv���Q��A���n5�5����79��QS��R��P����]��^��:M7|5�n�e�y�І��-�I#G��"Xf�ϓN ���ˣƈ���ج�)�����&IKH<��x�/�z�Ptz���yl휔6�*��eD�{p��i����q�D�����W��O0�����
�_�=}�ē�����W�E��4��'�T���9�;��z�B��O����t�t�&�-0�---�8�-%�E��/�^���V�=�̟>!�^n���&�o�ېus�q��5���,f��-z����k�ѥ�W57S���$�!!c�W[[����_��\l�j�����߆J����p|�ׯ�_���~����T�y����ӫV�Af����詅"䙨�Tq�g
�p08���=����[=>ь?��˝�=���:�{�$(,_=�wtV��KN��	�Q�@�����y�B��\\X�� ��h8��8�aR��		506>��BFC%��Ȋe�/6w�豿,�a�؅ �D@ 7nyR^1�<)��}��
`�ë6U�fN��ᗯ㔁�o��=�W�FR�XeI�<���bȵ�7Ð5f�����U)A��n�T❶��7h��V�b�V��En�!��޸�x�D�1aZ�S{J�,w7 �_������u���g����Lֳ�<l�L98� %����K��W����B��>"n�H����h�jE&��A��ޅF�J����C||| �����
G�i�Y望�l_��k�H��9���|ɛ��!i����u�:�'��8Ymmb�[['��O76��������!�h5�����>E*s��u2��N���+!A� ��a;977���S���܅Y-�׌V��z�`�����Fe�Ksм�V�4��f�VFI��]\H��ؘ�85�W��8�u.��E�Y���s��,7i�8V�r�H�	)y�G;c��x�ы9b����L� ���G�?3N����������R����7�^��9��N!U���/0usS��r2m���,��j�8@�5U��5J>�S�ӑE���Tr�4�D&c���Ʌ��s1���:�s7�%vJ�+Zp��u|i���
Lw; �5��M�1���:"?i��������'����}UcV�����	L��JL�{��P������ԃ�����Y@��P��@�t���ZS�Ư���)�� �P����l�g*W�%
ĝ�7��pˤ~~0͆۽�M՟C�����aʜ}��q�s���̺����_��8���cD�W�M��;3�1v�F�$A�W��M��c��dlm2�{+���=:��""�K�4���"D�����z��0����?�u����_�~Td�s�VAZ4��J�a�#��i����U���j�ϸGhT�W��9bOZ��"v�j�j#}��EZ]�R�q`��Ϸ��?�FO~7B���sl�@\�VO��F����(�̯7��2j����ָ�t�	���B
qtt��1���\e�����L�Sy��S��a�z��X��Ⱚ�_'"V�xTQ�!��E `�d�M��7'�'v��)�+�
H���d�����^��	��/����y�#�n�IOaq�8zp"Sf�(�٭�k�߰��A��*#��y�͔B����������8��C�J�[nQXY�ge[�
�aGG6��$�#�tX1��er�DS�����Rr���9�Y���V��Ǘ:8��WY� Q��+����N��hOrc��x����xو>%���D4
x�M��"E��(lBz
��5�s�d�I��MЫWha��,��55[�L�L"�3��K���S:�!!��C��{*���{"�֮nB/�����6�i���ݧ�k�)�����fr����m5~j�Qo�.U`J��Me�5�0�� �FW�F�J�1K?���]'�;�������'X���K�Ȉ̀���Ņ�O*�3�����9O ញ��nnn�p~���g��`��}f+F�з�]�Q��&_�����脖0F�]l�g�ER��?2M^�@��`o�[`�`a.E	"�1*���~T{�M"���U\f��EU�d�T{�"L��S�����lu=2<N�ᄈ6xM����G2�
<Ǣ���^���ڷAL�M���d��I��p��''���ZJzz?�������(����� �2��ҤS#K��0��H��?�=��i g��S{�Rgढ़�\엖c@�Ҵ��L�8�A���L�SF���D�K����!�6�_�TYb<��� ����a�-�4a3��0�#[�4��M���_8#���
D"���+�	l��:§O7���Z.�h�,�ɫFFř�������J� B�=�!��U2�9]\Vy,~*��44�YA�^bl�O�� ������#��r����di���.�K�ㇻ�
�J���(T{��*D��?17�}����l(��;�Q�[�܊i�Q]�<^�m?tx��ҳ�N\ۇ���$_�n��;q�QQVv��p��W��0 ZYX W����m얇��rOe2�
C��}��.#�A8s���9�i�(;��h�<t�Qy�7���
fJ�}"�����,��Z��)��M��N�:6<�i��O®�� ��Ɨ�/6٭ŵl���Έ�13�!�N�r���"��1A\�̛I��T��jc��O�YZ�0vg�?�;�y��T=�"����_"�Y� *P�O:� ��߽��ACz-.���SRD���p� ��XMN��_aRe#�2������%�n��jb*q����	�4��"�^�F#੧�]�E��斕�ިG�]���������'��Nj�G�����+�d(�s��pS˥��T�Y�����R����?Cdd���������<�ƿ�z����/�YM*H����G�-o�x�tsM�����a��}��!A\��Tj�YY� |s,yS�
ut��j�� uMM�s�ˍ1v������S�
�lx���|;�njJ��Ç�NGp?f|R����A������TK���C�=�eb��ǭ˖��������|��� O�*����:�R�	�&KX���%��f�GiSss%PTT�M�S�C���s~+1���u,��W �Ϻ��ர
����ո���b)�e�gߞ�#A���o$O�"-�������f�����{�!���$����2��q����G�l���?r%�郎LOGцhLφ^,Z�R�� ��������#���3toS����L�%\`���eܭ�����2M������J]�(���e̜I���Ϳ�y)	%9�*���!��2H����Ud�h���ݩr��	Y+/��J%��.TJc��D�6���Y�t��W�^�f�� ��nwm�UE���a����@�����
�$��ɉH��K,����!�Zcx�ml{�U騨�F�^m��+�]]��w� ?�T)�-�����g�ą�Y�#���0\f���ϣ�=e�k_v���,((Wbo��)e%�*��GL����qS����XT�*��V!� �{%��虛�%*%>I����L+8k]	�KLĪ�<h{C�M�+���j:�V2��*ON.�R�����}I	��r�==(��X�Wy��漂���P'd�)]�aN�|^!>�����Ʋ>�|(�y*'���ǹ����n	C��<�Q��(�
1�
OϽޯ6��ν�چ/�gl�)��Z�/:yA�$�v��݋���f���}kd2�'7�'W	�L�XN&�LQ��p�t��9�m5�X�N�,H%�?@�^r/jv�ٹ���W������6���7B��+S��i��W.=� @��f���}��qF*B�Ԍg�p��!�_*|��s��qHէu5d���Oʊ�14�̉3^����� #�s�Ou���*�(zY���9�xH^���x:-��q������tOKY:��Q  �yƨ�LO��8�%��/��N�k@��U���d�k�~�~<SSS��*sR�A5qG����\�mmf묵c�9[6�vY�.��?�}%Ώ�%DXL�a%��
�ިf,��J|%���]^N|�3P���/!���^�L�����T�U$i[���)%�_D���A?G?���dɪ��V�դ��'�r�}�P�\<�Y)�\?E�`�R��EA��@����i�B�^Q���q���B��5����X~��,��t���o.J[�Z��f�ו�����*�*�K�_k��	LNJzu�ՙ��>�P�/�4�^ϸ{,-3�Da䥷\>���
l�uY�_���'p��b_�Qaf*M㷻����I�!q�4k����f�֌ލ9%6���M5��n�Ŵ��޸3"&x�m���eo�n�����v���n�o(���J9Hp����D~kE��ЫĜ]��ѵ�x����A�F����>�U�`���g«�H%��[�)˞G'����)��k�@�CO����S8�ÿ�F�*���{Z�Q���-t���g�k�8IoL�eFa�������5�7s֖e%�,ɰ�#"uV��7%R]j��pb��^"N �S�E���{?����+�������O-2̘UV��<u4�����ŏ����Ã�:�Dj�����؛ɛ#yX_l>���p�����JIx����ȫS��K �����z^�6���<<�5.�dd�{��J���Ītx�!���K-����ay��sKKR��x�Il��NY���`�C.��Z��:[�R<ܢ�(�t�/e�Nݛ��CR�^I l�D�Ýp���z��O���e�H�rRbw�����"�B����)z��}� Q����*��<+562�5�LK�4����j].0��_)I1���k�`�j���"sSz�ƌ*���Xڂ�ɣ�%n#kV|���a?��,�qI���X�����**�)�Q�T�j�

�}ނ<؏�ﻔ5d/���0@���� J�\���q���\����,R�(��_>�$����m�9A@��}�iP,<\[[ۇ�v��#$���|)�6������i'ܖi8���ц��!�u�l��C�*��xg"�?�#8��>�_��>�/�N��z�o�-��5���O���Co��0�Z���JV$qt�ҒǦ���2�
�6ZV�jM 9	IϮ�n�Zu�uy �:E�(/����@�ze����ky��+��J�s|?���ĜGF�}���`��G� pNk�yt?�'E�v%��ʧp:��q
�{���(���i��-˝�|s�������� �S�rgy�*��<�k�NJ"d�^��Y7;gظ���`Wf���]f�&�Ȍ�C{���wC��2r�Cn�g��7ځ���#�.�l��,W�׽�d��Tizq��a�:
���#e++Z�\��
�urzgf�3�\��h�[cY���a���ee[I E�����!67���K��^n7���\����p��~@����"��3G1k���&\�0cȪ1}]�@ď�������O�V�g��F0��k�G1@�ɉ�k�%n�ځ"$J��D��)	
9̞���Ӷ��+e��w�R���t0lJ|V.� �@�^�KtW7]�'Ɖ�cM�]�V_��+��C����+!oDXRV��Fe�����&£_�o$�a��l*�q�&ff�n��Q=��=?��ʙ�Zb?K�.�[˻��Z/�"eJ�W��˅-�ֿ@�C�ϘI���;��E���Uu�����S��1�B*����_8��Y�a6L��o��!	(������"�R�:I��=s9�@ ���>kzfQC_�^���� ��
�߾�h(9�9��/�D���ND;�kyW��1r�9A8t"K��d�����sx�{���o���( [z qf�k���\�z�=����j�n2�n�k��"Ԍ��¬��L�����6�pz���Ğ���0L�W�n}�F�L�&KK��/����'&��vnV��<X9ދ� ���ٙ�Y�]m�ܣ���
�N�Ŝ��'~���  �1��N~d����4pJ�o��M*����܌eȩ8;�@~܋Mgg �
&���R�<�
)�
8������;	RF��?��~5�ئ!hj�����3o�RK�����0	��lQ���&[�k�Ӆ~������a�"\���u ޗG�������m���r��t�0��\�6Mޫ��Ǘ4�<Uzꝫg΂�����h��o�gn��ks���
��CpJ3I2ejtA�G7���0�0m��~����K.eUߋ��;��ρ�z�����*y_�˟o�#t�{�9�lrq�{�-˞�?���Dd% �fі��X��+�ɬ�������,ͫQ�=�+�',���ӧ�[��^>F���(�"u�4��T�Y��<^�~�~��zȴP��z_v�K�q<ڻox��y刳b�,�Q�S��J�9�K��W��DS���y)G���K�$|��sy9vfLq���dP`�'-n���o��@��?�aJ�xϚ' n��ނ��}���r�ϊ&7��=�ڝ��3�l'���ɘ�ͮ�4��9�jU٭w�ؒ#TH�;s� �pK�v�N��ۗ-�`:�ԍ�&b+���5-��� =*o����Ҁ���4�z�jb��LhD�8H��l��պ�{u��3�K!b,($�<Uf�s�(O燜��ǠV[�<�����qf�D�����.#3�x�\!>�Sg��Z��Oe;��[I��I��[�E��Dw0v3vR,lc�5���;{h�\�MȣKQ��H9�zxG4S����Z#�k{&��'�jnN���3����w##j�ǐ�3�J�m'��{4���c�~���c���؝]t����~�U��w���Q���ʧ���z���s%�r����{'^>�_D$�wd�;p�_��\2�]f��jo�Z�ӽq�>t9P�LBz�:�a� �Z�u���E�D��c��X���u�Ө߻���PvK�+�������'�C����wX�bT���_���WTk��\c�j"b�ӣ���"���ώ�o�������G��|��;��I�I� �2ӄD��j��@�9��-]�o�@����*]|���Fp�+������۴?��6DI��d�����N��gư���$����=�L3t{�޵6���*��~(8�0ppj�Nq�x�^�I�*�6JR\85�'��b�qe�xYT��f��b��*lA�]4K&�ε��� �ydS�zĝ1<��K���ӳ�r����B�[��e���4�"�_�L�R�ӼL�2�T��Xp���\�86��"-%���ψ-���Q�XJ�{kI@ ޷�)���������U��֙֏>b�*:��lU6�Û�<\\��_�T�Xj��ĭ_N.Mq��A�g݅�?O�%*)J�r@ ��<�
�E%	Dss3�@�*��v��E��`����I��\?t�+C���������� [,a�Wᯜ<0������Yvo�/��YZ^(jn6�"300(60c��y�t[�{x
 ���e5]�@a]��� }�H��E8�C�תhv���Ї��}mC�F����'ݖ�5Bhwxq��4�����L�
oM��5�����8II6U#�����h�B����ka���忯�¢~���/��3�t�p�Y%\:K� �(�Qf5dM��/����	�*�Cq:��K"��@��qe�##��e��E��bЈ���*�ŝy2}�J.q��28k�H��Ś���E����pP[����5�� 49[�WT�D���P�s����d���5v[P��yiB�5�7禷h�\c	�ߟQm���j̞����70/B<���>0o����s��`����{� x���x�j2�l��?:����i��S�I_�.d|�]󜮉N}1�l��G<��T�eڲ�Z"�媋I��"O[[[�9]�9�kqy!��)��JuqqQz��������sx��x𰝜�*(�`[�<�L����0L  ���#���b��(�����x)�]&c��v��dݠGa  6��)�� 0܂"a��D��zK�'�����b�����(0(ЖWG��a�m�"�v��ۢ�����iZ ����!<c�L�Ҳ��ITTG �h�f�� HJ=��	2)jgG�?�p�e��������t����;����-�h����{�6j.��@��ߏ��TxM���؁��Q���x�K(��׿��Qn���W\8�z���
���Gv�]�ݙd�x�����_�q�Ogc;ɶ�
�@(�}q�O�-����#�ycccy����I���>�ꢅ��� 3$����v�7����?���~L�}���_��R�E���o�<ݷ�P��,�c��	������icVz����Rh*UEj��ɲ��ru�FK���m��E�sl:�OT<�]K����N�z�҇1|�v�
�����2�%A�I�����o��<�fLUY;
{�g��w��,)N�}8��L�$-!)$�N� }����Q>�
,&bC��-C�w����+p[�s&A]�PZm�h�{`�䇒��w�'��$w_yJ��G��\Fk ���_Aty�/�(	�9)MNN��!�3�$ӈ�
�k�/�kw�����q�jj�aX/�����_5��1Rd�8�nu/�N��Ng�\Y��S�pq��	�t�#X����Bn䠣n����<��������4C;G���g�pW������ޣ3{����C���*�a�Gؒ���r(Y3�^ ���N�q� �bݶ�	 1��)O�R�-s��x�BҪ�v1��S�rΟ�Z����{�=aR&{C�,w�$��b�@��W�:`2�&�Ui=�v^K'���t��D�nh��oq��~a�,�%0#�=ȯ���l�f�%R	WV� �����wm���� �V���o]�p����E���P��ӋR����ANs��}�˿�L���;O���R��\0|Zh`EIy2m�v}�����<�<Ok' e���DA%�^g�1k�w��sY�7��c�,��Y�F�Q�xj������LLOGQ�<��	�_��]^�:����s_�� TU6�������!�A]�W�6����b���nlD4���bem��M�/3*N_�2(nm%<����Π�읝ZB�/Eݟ�Q^#�l����E ���ظ���-�� V$l��:stH��o׀��Ş�����>|H�a���-)o7�t�X��߆��k��䪳v�MK��y��iz�zT6W�>�+i����8��_}RWQQQ��7�S���(�c<�V�0�W��2p��.�#���=J�?f�qס����Q)���+�?W�'9D�q���>��y��n�{6�X)���u_oS}��է���o�	_}��2aWq����Xb�(��2�4%s�N}��)���y�ξ��=���w�����6<�����ȵ�����E�](�M�L�&.S4��r��Pc#BY������7p�6�~(}�b��8ѐ)���j����O!�?�@Ĕ�Pq�8wd����Z�y1�|V�׸���� @�c<�fQ��|��Iߍr��g��2�u��ss�ʩa��h��F�_4����fZon���++(,�����+� *�B�ɜĒO��F�r[`�2W�KnB��$��7��N+����K+���,.2���\5�.��EΑ(6������%�x�]���v�lNۈ �0�� �<$d�\���D��qu��g��5�ο�r,���e)��T�p��E��E���Ce��������}�+�P�<\NF!���g��[VV�3w%_��e5��1��]v��*lc���	W�A�rÒ�m�Bbϫ��]�L?�oA� ��%���)I�i*9j�G�,���d�]H��O����RI�o
�Bfm���L��諸� �Y��P�>%n���=���	����h'�A�3&��������B��"�X���F�Y�nD�	���Txx�C���Y�H�����]�ؘ\L&�5`��������L��l��K��2�դ�S�m�̭�[�saOdz�Nn
?�m���~��_ۄ=��/ó���y	N�V�僆�t��<�R��}��|�U߈���=��y_���%�b�exÿ}���%�F28T�Gb���GCKK�;����B�	�ͽO9����y��׿S
����u����Li"�l7��X��Bp�p�LK��z^t�����M�g��cTUU�d2��+^T��d��`���[�^�V�@���;����fBdݵ�#���]'Xhh�B�����[���ʿZ!u��֬_:��=�ǰ�]�����=�Ü3�˧z��S��&f戮�כ���4?7XXad[ ���3[ΰk첃���o#�s3�V~����K �� ̰�-7��߽3����U���Q��Q�M�Α[�������W2<3�p	 <��\�ڦv�=���J"�Ė��ggg�?'
=���qpT���6;��7��V���q�F>P�q�j�h��#TA[H����-�kS%!|u<�+�����K'�'�^<�^��]���.M�-�zQH%�A����J��m��vv؄4�s��c�bb�0����1#1���0�i+3��i�����e�s���[
���Gg��x�
S�^�Ih���bnm��+$�V�6*��k��Q���j�p��;9KEYS��AQۃ��� e�ǃA^�1��1��	��l��A���m��q;;ِ���8�
��#k��%�,�S��~�U�wiQ�ﱼ�y{�����1``�	�K��B� h��޲��M:偂Ґ<�q��s��Ve�1�!$^(��za�*�[��}6옒u��u`x����3���"��L4T���23�bQ��o#�HH�l|�H������m��)����N���K1X1�����Ҳ�>76�� �
ɕ���K��ţ��n�a!~�3?=�9<Ԃ�$�:�[]ڇ���"�G���^��TTUE�)K����pjgn�y{�v�FݟvKw2���3#�:����ϖԿ�C%`"[��=_#K��덐%�1�$�X\�i6S�=� 426.i�k���`>��9Y�{&���MG%�J2�ֺp|�~����q"��B�l��/�Z�#�I�}.o�4�qsu�SO �s2�b���		�j�]*֛rz	�cĶC���5��Þaba�sG�լ&%C���ȑ��Ĥg�D�O@�����`�����D�J��  X�����]��~��R!�ks�����R݄��5�c� h���!���x�������&ؘ���=�E3����:�DsY[��]�P���T��{��ٙ���U�V(�0��ǉ�reKt�C�H c���0A�5)�e;�n�̢����{$�!*�_��~�Ժ�'���ag/!��',�ϳ{�l)C�(M�ԣlq���Yk��Q��qߨ�a�UJ�&�$-=�DT�"�ט����W�C�8J�h�#2F����tZ+�$��j�k���VNz���ܰ�jbh��H�2h��-'k`hT�d0�v���ċZ��`5��&�t㫼/��8��O>rُ������4?ԉRhY���3��n;nL�u͗�S3�c�_$0���O��Z+ؐ�r��2ǟ w��������r�am,1�>��2��aQ�W]U����Q��,��0Ԭ�F����׾�"wN��=I_�UgΙ������5�w�N�K��nKB�A�d1s��ZClI%�N�3_�ՒO��^��;�┕�W��B��~�fo�
�Ah�O3UYx�Z��2�&?RW����  Q��$ë���51au�C@�6�׊�hIh8�Î�R�W�x�Bӎ�<$`ec�0��<i��3��4Gw�=*
��)�l>�G5���#��cJO)ss����EJ[[[_��g%�Al�x��}e�T�`�:{��r��gg�**Tz�J�[%�4S����Cu�:VT���&�{�z��1/�_�7o�|%��R�Ğ��P�ؙg�lcj�cMU9�/I��g��0��^����P=�⁬m��YR�k�T��D��w�W���	2Ǭ�]��L�6#��))�&*E�ǫE ��L�  ��������eM�zT`��#�/g����^؂W�,��(Y�ٽ�֖� Y���~<���`���++V���6�4P� �g�e�H�S%n'����V�n�XXX���*B�c�����H�-к]�]dHH��e�ʕ�
�m�W�WMDXCs=W}�Uh��y3����{�� ��S�� ��;_pz���$��/1�8�Ê!:���B~��OH��6���L�B�̾��CG<��e�^2��aف��l�p\R���I��3��Pկ4�"#!#�aOwvv���yѩY���"=�ݸ�V��	���ٱ�4|��M�`����U,!/�Qr��J�٦����	j#��F��)'w���s���h����h�HmKK,�`FΠ�lh(��nqWd�p/��,�ܙ��`����d~�BY�����	뼊����r1��~��F=G攡s�Qh7�˗/w?�Ж
�~�~�a������A)�z��h��(��H��4Ғ
ҥt#��"!q�!q���4r"u- � GJ#͑G7�o������-���;�<���3��a�,Yp-����(�TèioϨ��??�VW�W%�S���^h7�}��F��E*�C �%�k��(++300<~@����/�p��֏M�kB���C&~^��v���i�=�866v��I$|xZyj
��@4˩��Xx�RË�����kL������"�i��>�jjj�w&� _Z���b�h��t@2����D�]O�A�銶���q�y�������,@g�:���`��g�e@$.'��>		��a�����(�U��k �r}�'�ӯ�a35�"3 )	�)�J_?�R�;�z~}�U��&��ys�Y]��i�1�[uh�OU�pI��OՋ�����d�BU��}y�&���^픞�b���^x��@x��E�A�2�-�CvSt�&g��3�8$��'�a��KАih�����n�i�[_�X��#��i��>����<j57���t`q��Y�����E��_�c����'Jƫ�9���[>�d�����Ƞ��QB}_*bY��I��1��<+;e�e��8�6�`r99﹗�۳.)J�Ę�klo��Q�#�O�m�O��:ï����WjU1�p��Sb�}��גY<Z~��R��� ���w-��}6�i仞��(A�o��߃��Y����N�	�e�P��i�s[j�WҴ����a����T4$� ��7�Ǝ��.�����/;/����U0=�i>��fa�)ħ6���0i��T��������\�:�E��E#<��%bVup�i�}���	�P��@DF��Ť��ߓz��z(A�����L��6�.�>Z����������`���yO��rQө^�i��{�^~��*�w�gv��U5�-�a�K��Yţ���D^�"|����L�QK��_>�
�?��3j�aM2U*a99w�t�B`AB�!_Wʶ�2�ո<6���<VT�S��������A������b�\%y�}�����%�]���;�_���iĴ�����R��N��r��5.��+B�i�0j^�������0��Z�dEvY^�RLi��I��.�-o����O����2_�\����.Տ7�,h�@8ɜ�9��p�R�w�t�����(�������`.�lw�� 7%5CY�O�
~pxo�3��GY �hoo߽4q�im;]}��ӣ�,Q�-h���~������2��_����w�kF��;=����>t��U ���;���.:2$��/�Y3����xݶJ��G�a}�E���̠Kb�)u��$2j
I�d�9)��79���������'�-0���gѼ�p�yI�ʻy�9��3K��nܘ��g��{��%pu�-�a�V�P��zXߔL�|���ǝт]^�L���\�:ڔ8<wf`bS�(�)\�W�!��S���\��P�ٱyq��/��]ؿѓ�lm���#aEE4y>��{��h�??BL(���>�}Nb������i���ی6�7��d%E�y���bT�N#���;V<ɜT�VFƮ�Ο��2|����:$�ڍ�w7���vF�r�wrܺ�SPA�(�j�d���#p{k62�"�W�f��WG�)B��qc`�f1�jk�3�iS���,��VQ\�`�����ijfVn�=��;Q/�{L�@��},u=pp)�/��}�=�'(�U�"�/N�'��@F �+��� f?$��(���{<�P�X@����66@Mw���f%  ��LBº�17왺�
���+Zb.*v�۪�%��]���<a
K�	#˓2��bA>)��0��o��,_��>�#�� �u+���D���IɅ�{S��m٣i����kj`��QQQ�[�XV
GZ�%Yh�y�ȥ���/������-�W��&��������]�L�+�m�[b�2P�VcÏf��Jw'�O�hh�dC��������������N�b�+�99�6)�\� �� 5v..�6�H:x�m�J8x��3 ��q��+6���3��oi76eޜ��#�����\�n1Tؒ&��ݗ�C�T�g�)ι���ك��+���C])���#�S�a�h�w����"�u����l�ӪrP0aq�V�����������q�'��n`c ������{h�C����͎��P�2�M����{��6��ty���R}g{]���%�����wy�D1f|s�lvV�ӡ k���гf����i������_Z^����S�����L.�����C���՞��+R�r�`jx�h]�D�D'*=�ܱٶ�U/'�m]�P��!���_n0)^�<�7�����Ћ����!8�����Խ��\\`Q�ar�\���Dh���T-Z9��������ͣݳ p�(���F[J5I��.��*/�{_���D���i��~���~�A������q�7�־��Y�]�]���M���^��n`�=����ߠ�:|y7<�CC.L��.z��`Uؔ��[a�k�yl9���ɷ��y���L	6���q��ݟ.���p���u�ȍ=���o�Uz�j�8��P��K��Ɨz��	*#K��3�2�����ڥR���{=\Tǵ���.��%����&�]��;��]�H�L����}V>[:�T�z�zz�ր�v���z^Ry�"d�0�2���eVU(��F4iU��-�0K>�� �yQ[m�{�Kl�ר��P}��1@�m�I�Ν;)��/P0���%5��ߎT�R�Ce878���Aa�>A޴�7h�B��g� 4}�uc�s"ڄaV���Q71 <卼�U�5��7����p�C��0*�8�@��2|�E,7�+ng����]�[���G���i�_k��]�!�;�: �>Kr:$���ȉdף��M�U$0�6㘣�|eb���3`!(�#�p#}���<�q�7qR�1�(!��g���ڕ=N��Ļ�9���h]t�X�t���XV�������q@#��O@�5;�U����TG )�^^Cf��ո�$P�'����U�ʟW5�/�g�d�J��7`Tѝ�]�nO�q�����7�p�ҘR�E�`�; R0�R�����J�G3��`�3�]"�j�c[C��ef�H�%`O.���Kf�0E�aH0[��+zM�a���!~uXXXBO���^��r��3�7H���yh�3��b��x�r����s���r��qF���ŊP�����$�;x�S�$xE�|���t���`�}m*���yb�|���5�w�mc�?�<������QԦx�R[e��I���ID[���fm�K�xs��Oj\�RB�F]6����`O!�����T��b.�poh���)=y��w�����@�=��f)���'��	�l��)Rg�h������y��_!��ng��[Qf�w��|�I||˾h^^���H�a���aA��k��Ak���GEA����2�J�rP���TV>]�<ɫ���'z�+_xye5�KQ����Z�A2Q�vq,�p ��\l��?]�(~WW�`�˓��oCJ��i�F��r��U�}��R�ϊh�����>�["%aK�ic=�'��	��IF�^���{3��$��I�I'F�|�o��KŘ��������X0�x���~@|r+���Ј.էf1�z�lhu��e7h	�"��b��w>㊜|�m��%�?;���ۡ?BR�	={�5(X��.���w��";'(���I�w�fv
#��t~?t$oce!>>>���^�xkV���T3ytx����0a(��� ��ߌ��,l��g���AI(����aOU���s��II�)>���������J|i��6)R�ػO^	�={4}ӫ����Nn�L-���=�_���ٽɗ�(������}�og��1B���,?��$w��yy	���$
����2�$4�kǗZ�~;�ܤ`W��V�Qб*�A�/<���`|-��˜��=	�a �l�U�%���T!�p�U�?d5405��s_��\�����t�����6Z�/�YB�8H�N�ɽ���$7����^/^�R?�~�狼���}��)���>�ӹ�x��%)P���j�4@�c��|@�zG[(����3�O�Թ�����J�+i�iC����mpvsK9��<ޫ=�Ƅ�>����O�l�̾���9����O�*��r5��*�>4:�v��'�����
p(�Oe����B�q��v���y�%rz�;�b��������(���$ã4�"���=��B��[X	Ѣ�#
=	�~�݁�9V��!����<3^�ێ��&�1��:D����ѹ
[�]Q����x{R��E��Ɠ�+ �J�2����/�d:��Ƿ��T������/������4�K�8
�
���` �4K�K�]Yْ1�yԶ�e?Z��W�g�X��V(L�G'S6�=bN����b,x��Sz��y�F�M�rٴ�uu�)nkS~~>��8��BwO����lA��z�qr÷9��G�����+P�K�+���sOy���l��6��+�a6$���c�\�����;�!v	b�Z|�Cy4]Yƫۡ5F2NUwt���7o9�@��'sz�|"�W�ߡAvGj�55Y�"t��^9�YĤIHIJ�rÿ(OMI�`�_9�<e�V���!I$�7�II����ͪ����'����Ձ1~1����ZYp����J�$�����!����߽p���y`g���<��Wa�4�_�����Q��@���,a,}4孖�o�+u�ϖ~�ƫ?��H��僓���I�k��)��H$���a����)9#������J��G���0XaQѓ'OB�f3X�Ǯ݆;�����>l��}b���[U�Tն�w��}yy�\ތ�U>�Ȉ���>�ee k�%y\Wxq\��l/�����0t[O�����y������mn�nK�B3�_�`2����iH��	;d���2���xx�|��#�,�<cp}J�d��x�z�����\b}B��y�7ho���D�g?;�cM�E2�2���q���ꥥ�;�'ja�p�������/�W���dS�!D2��ޖ�@"�����@~�?�gg���f5���N*���ۺxivy�$���~.����SG�/��E�:����-�ͯ���o�NVML�/l PLtѳ����������Dڛ�&K)���?�8��H5ˊ����*��mA6|�: ��fr���}�l`Z���V>I%�j�W�eI2��U�����z^^������kR^HP�ǒ���leO�p���w{�P�ME��//���qr�J�;}YS��XP�$�p�]�/�>󣡧��@�ɡ�c����������=˻�x3�8΄�qt�)����Y)�}���_�~���I	No��B��B�d���O;O��)������xt@`�;;�.���V֕������B���_%�Χ�ں��.������R��,%Q��uuf���1V2��#8 �z]����3큁%K��������@Ve%eRR�eǤ�
}3[�>W3/@�Khy���(LnG�����@/��g(/� o�Y,:�Kn�+�ܹPw
j���Ow��~<��frBf��ez߲zA�(Ԣ�5 {��������L}xx�?=+	�)#X/��V�MIC��i�9�3�>�<;��:�A�$�!99~c���h��bj��o�����2��J��L�|��4��	�ckr%R-jK���&��9Y��3�M��M��_�s #������`]�z�8��CJ^:!ީ�}l��~p�'  j,:�z,�j��8�~3;��p��[3�ǘ�YA���;��&NG�T ��{�=h��qyy9���穥��`���w�3��B`���籛��NZ��$uV�܎���i�"�� QW'���(���E΢��&�R�:L3#����^�L~��=% �s?�Q^�p��p/n���\KG^�T}!I�А�[��e��b$o펏pd{�b"炋^��u� i�q	r�Gf�Mdk�oC��5�<��B�eYss��wq����k�B/��p�'㫇���N��}�f��!UnB��鿣�Bn�%k��R��a�u����m`M�� �����ĕ?�p���ol���"�'i*���yXg�wm�����.D'�Jq�w,��:.LR��B����Rw����`u��U��<����p Xq�-��7��1�N�sspR��4p�4s$^��%���B��K9�&~;=���p��K\L>[���
��I� >(��C���nj�X��		�e�.�kl��-�>-��Sn�=/CUʺ��o���_���LJ�N"f��yR��'����}�I����Iޢ�^���Ѭ��7�]��._�XK�_Me+J�Y(�!>Acj�΢����7��=*H��83g� ��*( st��0�<#{̌���r?�c,}��]j}�n�����$�F���5
�1�(]��S�M�2=��~ ����w�~��Z�	��ι0W�����K��Ϲ�m� ں�E���e%�3�	�M��إ~T�,��z��A��N����,�}�5v�C�B)�MڛF��u[,�V�~*�y�����G�����7ط��׺��7M?B��o��Ǜqk�L#�f9;&��&=#5�K5,\[�f��iJ�v����c$JF��f�&���;YmgG�Am�n��������.��A� �ˤ�]�5Ts3�ɮ�L7]�tٔW��ۀ<�I�	;]�"E�.�|յ�"� ����ȧ���𜣃 w�k(lmm�ӵx�Tr�hk��NW��ST����4����>���2}�p�G`;�C�l��Wƺ�6��[������P^��tI+���=�����4ݑO�������(u4����بR{� @�Y�R�Ǐ��3]c����TTU���9�4�'���?(/�M<D�ޱ]Z`�ؘ1I���{z�I�$+K6d��]������*]]x��/�4r��3J�b���F��5�"�P���0ꤩ؅t&�\��;B���H'��l 	''����~�<��@~���q1@��9�e���2U���ID��M�_��X�~���hH�1H�6��<O�f��}[��mb���@=ʺ�.���@�[��X���i\���˙[XQA~�X���^;M�
�V�[��O���lq`��3L����v{Ln����H�'�ʪ�M��]=�zJ�[?����>���5�5E5��>.;�JT�}��L�b�wd�:����ݰ[�C~��/��C�|Ίi��η������L�R��p��]1}e�A$"�L�>x���%''َ���`,J�2*l�!
���3�d��Xs�@1k������M�'n��~�,�A�8x�RL��!��$��'K�g=��|nO\�����`�dt8���h�I��|��/�Y����U�_���h-�_'zh�9!�D��r��u���1����ؽ�oPA_YVC#�\�}�P�_��P�u�~eR����p�c\jSx�,75[j��9c�'������6Ud�n��K^�eec[z\�3�Q�9��=I�C�q=��#/��q/v�����uw�e��hѓQ ��Ȍ�e�I�[�J�>k^�E�]��2H����X���#�Xkn\����<EVNr�Ow���W�{#~:V�y�xվd��D,������X��95uFR���yzhv��Ƴ4�%�W)QVV���pk�w�T�(�]{���o�;y΢f^>����
��0/��^�ܡ-��xy�b������F�k���i>}����iC�5/��#8ڙ�A�"Y�����	N�J��R����y����^\V�#���K ����|�ߞ�em�h���g�y��L���N�e]�æ���C?��/�_�IS�/�G�H-+Lg+��RQ~���d�/�@��`���1�Wao,-%�-���%�(m[�F�D�oyK�@)���o��%$g�c���~�A�pv�,�S9�4Rk�Ixl �	P�1+utu�3�T:��m8c��f�F`
�*��O:���/+�F!��	w��e�����纽���~�ዋ�����p�h��v��G|�h�qt�^����|�uTu�H�`R�rR��̬�U���o� �6�W�w�7�c�#.qp��_�9��8��554Sj�W�1�o�p�ؕ]�N�e��Z}�.}j>@�GAFֲs�).D���r�5��_w�'�
����CA�3?1d+�i3Ew���T�JKKG��{���i���������{C�Ѿ�@�ܜ���+z��@�)�k��V7-$x�f�ô��WœQ,�g����7&��p1�ݥ"70r�`�h�C"j#y-!I�/�����/w��y���J�!_�<>&�n{�|)��+n՝Ķ-�MR�	<G��:�>/p�X�n���8D��E��ӭ���V_#n�� ��Ňm��.��ػ6;���mGGG(���Æ���ӫ}������E���O��zp�!�������G�t¼"�C��g��x��k�n�쫜tIA?�`��jt�ך���cg ��T_��8�Z�[.z�'�$ԓ�5��;ͧ��K�����{��m���>V��-�쵥)I�5�j���K;>�����~$&�)�!���R���27�<bnS1Z�^0�MK��jDa���/��tQ���͟����$�-�/�=��o���)4�`�,D�C3ø��h���޿m��c`u[���	����z��(�o�ƍQC����XfLj�4�&�]2r������\��Q$�/&�dzv��k4��>�>}?�n����>K+���f8D����0B<w�զ���J�:8`�1�cz�
�|�_c�*�����6��g���������QWf	`K��Rߥ�5-)O��[�an`���͐=9=���u��Y3�]k��+���@��V���G�U�eq������UD5�yQն���l,+�0�2	v>c�u
-���!�ŀF��Q#ւ�k���,,<� �e�}�̎n�9_��߬ �N&L��c+04������%O��<���-M/�0զe�s�I�ehH�[���X�l�^��kk�Kgf�FS�)}p]."����&�ۇ��dU�#L]���W���%5��'-��5k��V����^A��	�G�a��WL�h��pu�Q'Q��p�?׹���i��F�^e����^ߋ����x��������r,�W�ixV�>O��,,h-��LN�B�d�
		�@��!8�t8j��'Q9�jEu�1�({nE�E�W��``����&K�����=2�g���9m�7���Ц�yLK���g�=���oLg�A!��̢��~�X���6�#� ����~�.�WfY��V��D��񾆣�wd�,�����)�����Ƃ�a�{w�{r_���V�4����_k��#��Џ�x�|��J���OH���G �E�2:��zs�t����y���9���h_0?B@H���F�W�~���ZP�B{�VK��#y��8(�?Pv|�l��
����o����"�:�}�g�x�|�5���0�݅T�ّz�4s��Z�=�L�9�R�,�j%��-�������¾U�@�����]���P���*gF_)�_��g�ma&=��5�1{��j��!�#`�(�Z%9٭����xYb!###a�e>����p��ϑ�ڸ�
��B>�d���i�
���N��!YQZ�Da��J�7�r��V����vM�C9�'�hσb�����ud��v%T�A�">ta�Nʶ���Jh�����I��=���5+�9�|���"П5���
�-�	�5C�����J�/��R��ͦQ&��#�L��P��l�"qɉ3�{,\��%��J4_���.�䐈q�SU.�T��a���n���?��ոB�����˽��n�7��F�e���{آ���O�;s�.%^�]��8S��Le�Yr�A�T�Ε��YS%t�~뒷�t��6v�}��{LCi��("�"���nuվ�7C��~��������S���V��-I�&�4����ӆb�����A�u�Ժ��?�'߬mpQ֕Z��G�	Knll(ɮ�hh�PFO�n�9�.6W�/&�h� .{��tsqRxF�{��:�/��7���n���53*K����+5
p$�����
���md�hh`��/��'q���'zY=Y=�j?N�
�{]��M�PWJ����T�/� �%77��m���K�*����Z �����{Ve%�g-��UP1(�]_W�/��x��s9=�!!Uqq�o۞kE��������O�
I�ؿ%�m}���G"&�Ód�A>�h8�(���L�Onq_J�1�u05e�H\<>l�_Գ���;�AZ9�L�.�l,�\���@aa�R�w��ky��?��53_�ǥJ���|6����k���w�4?����M��J~�6^TV�/Sʧ��8"�b:]Zܫwb��_��Lk����F1�2��3h�Ŧ����M)��&&ġ7)8�}��ρ���\{y#�N��zzz��p���� �5��+�`4������=�+(D�a"/������N�S%_v��Y�_��gW�*��I�r�T�846�[�40�t� w��\�L���z���s�������a�!��F��c]��R♖�k�S�e5 �/�;2�]�x1�?,�8��Bi��SG��Ϟ���z�?M�櫫�µ�ͣ�Tq���×�r��-�%K���
u0���Y|&7���A�VE�����AlJz�����>8;S!gK��V_߻�v����,�.���ߋ8���l'�߆|�o�uQ���<b�Lv�Q.<p68H	�	�(�S��� ����������c/hѲ��A����o��6m�5��p��O��X�-�5��ٰ���c��.���������?�7pV�u\�}5�Ak��i��UAm���
���@�q�2M��ov"�Y���)���P���j��Nb�B���+<1���c��a2+�4�EgH3"�d�n;����W�fۨ}�*̤<F)��b?���j�7�Q`f����ԓo$B�����ܼ5(��h�L�-𭯀 ��7�C�/�$7]�&]��de�n�_'^�H�Vt��������1)Z2��8޹�2�1�T�����	��y5���/��\���/|����}��(�'�Dv�4n�����`�b����20��8"##���/h]��Uݴ��so�)g�c�z�'���@->�M	�OK��^n�a�Q}u�����/����ti<�l��42�܇ް���4Sx��Ih�����2>&�Ǩ���<[+l��w��υ�8��.�R�z������E�A�d#cV&���|�~��s�;���y�QK8*��$�/�Զ/<��{�'���{)�|;����^���946�.;��W�U]bx����R!;X��6j���X�w]��X���DO�K��un6}�Ì��ޓY��goog��y����MƗ����}��+]����Iϊ��_�bW���D�������R�[__&���g�L���G	Lg�,�W������N�ސ�312^�e��R�س�����Ѧ&|�od-@ۚ���Wkq܏a��6^O�zO��\�@���>ё�= �����M�J�U1�z���lh>\eP\�S���߿?���{M�U�_�9�9��
����#��h�U����ؐ�k����_#�>;�C�O��_ƾ��FM����UoF�t*�ҔtD��Ds��UI���,��+%�E��g�i�wl��>�"(u��n���~:��)�C�}Σ����oX�J�r��E�?3,,��^R{5BC6����^%��gˠ���D�>R �ce�2�R��r}�j#P���vg�s��)�����'Z��Mz���
x���r>�ׇ�i��	��S�ӫWv�`
棣��=4��=�?M?>AA�ׯEI��j�&������?�~C�NU���'�7����e:I���y��z�e,�nȉ�K?=͏��.5nڢ<�$��-���w��'�.�4v:"n�Y�E?e;鰍_j��Z6�0�'��S�LK7�Y����CNl����;���.��;�}��`��|�'����������O7ԙu0�E���;�Я��К��濱����hK���M��KnY!�w�7�d���6������ލt"Ź�],�����~d�q�_�!�k�F��=��8#��:갸����xq!b|��G&�S�|)ݭY}C]h|��c��s��w���]�T�^{G���Y�20��~�ĭ��b�(-U�S�d����!I����%g@��G|q��3��ԇ��6!T�'܁�d18#S�a�Q�H־����`o�*׿�# S���R;��=�6}�@U��ڨ���ֳ�6_���*����;��������x���]ߏ!��u֟.�E衸ϻC`E]檵�jY+"^����|1UB���h�6���H�ɬ�z%,�<9��i���x���[�bc|��F�_�U�D;U��S��C��z����Z>R���U[1p�%�N���a_�PQ���
�괉�jl���"7%	�P�X,4&..��^sTh;V¼ �Am�Q�"�G#����y.��*v��B�Mo#ȿ){�?����zj��͐�lW�g�!ӗ]�*�r��y.B�����bM�����0v��ޚ�T�ۺ���@H��}��EA0�@f�e���pX���N��c��=�H������ʟH-��9��wy�Q�!��ԝ�O����l�����=����]tuس����Kd�G�`]���իW|������ʭMM�G�i�u�����G����KM�L'Y��;9���|1%k��ì.�������mU�vG�"�ݹe�EH�D�L{��(����l��:�G���:N�>��sN@�GX�bBl(qf�O�*�K�'0C2�`��T:��	����7o���A9��k^+�ppR@|w��� D�
���]�Nl�ӗ,��S�w�Wj��'[`A"�f2kD����h��˰�a1���ɏYS���_>�d�%,N���	��ϳ���Mֺ�{��q�bJy-k}a!b5�G��m
u2�e�dr�	k��,��`��/o�^��R�R?�ص�m�Q�W$���Ӓ��II��:������v��.�yd�}c��9T'�ދ8����s�7�pᲣ�a���J����ڋ�?�h�,��U�Ne�O���ߓ9��R:�<D�b�4��/��2�չ�o���@�B�L�ON�V�_�Ũ��t�����ա���RP�ɏ�COnf<=�0���B��ԟͷ���j���R��0e���x��]Y�#]��7�����ďӚ���ӭoa9��.��Tw��Đ�|�2+/����m�zE�11��$q�q����Yi2$1pt��E��ꪬIz�=�4'�����Q�'�kDE��NU-~:�a�r�rZ��X̚��y���)�-٤�,���M�\?�+������H������O�q�s�Lg���rc�R�e�����Z魑]��T��4~ Lɩ���DL,���1hɽ�ND��țj�aO��]�I$�W��A�>��;�Tn)�p���ݩ"�ʤ��-=V=JL�մ��JJ_��S����̶6�c�=U%���K7�x�ُ��O8F!�9_*�S\�����e�#�C����`Q9j?��ݚ��Z���Z�<^���B���S��QH1& 
%���Ϋ['���򲙂:�b>��MM�����<Н.�L��-,sᗛW��7 ��p	8;_�`2=�v9n���;[m'�`�����m�_. 0�5���A��4�e0���pt-��2�C&K���	����k%��z�`��;'��	��I񲌝��i�~���8�\]U���=\���h�g*!FD
��w5萱T��5X�qv�?ޗ�<"��u�B��Wk�,,b�$bB��>�JJ��z��$��Y[ �q��|�}��#�{z�5V��p���n;E�
��AG%(�UCC��8������=B��S��H�ڬ�Y�K��}|W���Y,+y�N߇��c;i���eX��[9^b����~J�og�u�|�����:��L�$P$tcrr�TJ��_�H��v܊z �~x��#$i�8�c�R�(R�W�����A���6	��48Uai>�����|�Tlt,�|U7C*R��j�Ӊ��Q0Y�n�R�Y��AmɳUC󈰽��BEy
�����<7�.�&�lx~�	9@"���	s<����uʼ��Nb&��A�KAÏ&/^�|;%E����CS�$�i�Q�d���3�Kⷼ��H�}͕n��G�MR�u`�l��suuM�e\K�N��^QI5�t���]k���~���ܶ4�̞)�<�&ű��hVFWV��}�I�Q��5��ܬ_x
"��R9�u����I�Gw��~Ŭ�&�E���?�7,r�}���)`�!T�����������zP3E�q�����Y/cd����ѱ���U�Չw�R�0�꬚�PG�~1�35�	�?������|?��-(���dv -+/��[`cs3�0OWG+�����b��r����B[UP=KP��)]���^�[=�4�rJ�	�~1u����������P�Z�Ҡu�d�/U䇷�9�`�I�^��oR�����9i�<x����.�'����.b�%ߨ��.kk���_T�e�M���:9�r�f�G$�t�NNN�\��/<�|$��RE���n��+5XZZ��X^�� n/S�S��\�X��^L``���O��̻�/�P�fǿ�	�o��Q^%��d��$Ϳ{U)2M%����خqESf##U��^{~��R����Ň1q19%%�R��:�_���e�����GQٔ���}�o�c)y�Of�o/�JI����Tɨ��-r8�ΰdsOo���)�!_[�3[.����u��EM�NyUTHu�R���GX���wf�%�&詯�
��=�?�=�<��6�Be�A5I�{��'T{"�:4���,N:��c�iHd�Frh���u狉M�)ʎ<�H�zw�9�n3?'�I^�O��J8Vf-���VX��Y;]����/C'�!���p�3M����D���+_o�塼r���D/D�G����2]m��D�58�����Ðw��_L�n_�`�b���3��"]��&��!�������4Qg_k^H-?Vs<���j�z�,�&$�d��Yp]ݤ��� V\yz*���RN叕,5����-�v�T��E⬪�ٸn���j��#��-�j�/4K��`g�_f_�Qc����T�u0� �2�����I/�ѳ�����FR�=yr�5`���r_3V�H|鷉u>�s�1ͼ��E��_�qK��68��X�\'jfv�u���IJ���m���Nt^QqE�e�#��V��쐓�@3��N�K��ѴR��t�P�n��E���$.%:]����xob�!��F]�bs�&z�R��SG���k��"d7���h�h){��f�}��tf;;;_�n�5�f.?����phIg��%�������wN1�}��fYV�_�T�#Q19
�(���+�h	��xE�'��#�.Ɗ[aXv8��Vo�qˮo������
�Z ^1 �>����U
-'B;��ϰ�݊7� ��9�s��D���H��-X�H���:�VU�g�(#���L�5:S4�_(͔�iq�PR3j�Q����?P|�߉�4�fL(>�У�ye��qKӈ�ܩ��6��g�,��m�i������'�����{r�Ҕ����'<�ѯ�@d䴠� VBk����IZ�-ʒ���'E�_��t*w�{1ܹC�7��u�@�L��F8 .Q�����W����r6}O7){� ��/��+���4./�����;� %D�|��%��v���0/��<�����Տ�S�`���޺2�LoW�7�*��W
JF�84;���C_��b��u�	����/�5~J:al�wb�,�4��b7�ʟ�����כ/�T�����������?��W}�s�]3�Q�|}�|������OO��Þ ��ޔM�<Dmx�{�˧F��qh���J�b��v/f�}�y�`�k<����૪�K���y4������酔c� ���$�\��ڷ��7>��K2{@�vzE�ճ�<7�g��x ,0�ƅ�����4�	�wTf)=�Ru#a6��C|� p�B����;C�4���[f�:��͑۫��h%x N{u�j� @���R,_�~�u��i����A�|���^}�{m�U�?�0�L�����M��oH���	�p`�z�4Gl����O���۳�/�=Kx�n&�����֤h�I�`ui8���G��I͟h�
Ň_w췰��;��n���b��/h���{H�[XR�T�u�H��������|T V�6ҿ�5��]2����K���d�����m��/;�< ��k�vNHP���P+�Co����777g���I.E�NO�`�D�	��÷\�$��vT��Ȕ;;KC���m]n�� ���j
�$�W>Ϳ���{��A{�5 �T[��F�?=|`����t�m$!;"ćܪlhWf��垵��ڨ}M��R�e����	����I9�U8:E�*fScg��ޜ�bˍ��gڠ> 3�w���u����[9B^^4�r����[U�3|�ᕾ�c��賨g�.*��g���5p���KL�sf+�>(�J=�,x��tk~��I��)9���ن�T�!%ؘ���B�V�����h����p��H0c�3�X3���흌5(�E������u���\��n�����K]�Pt�fD��)�K_�a}�a�s�
�&bO��x�i�yߣ��h��k��7�SX�Q�=�������8�ĸ��1��qQv�ք���4HHJw�����t
H�Н"]"� 0��Hw� �t�0 ����{���/�s�s��g�}�Y��1��\�_M���c�R�./�m�\!��<1i�8�m�b���SK��OQ�3�y�Zt�U�I����@b�ĳ!؈��N�����I/;K��A!�<�O6&3�`h�� *� ��=�wi+D({R6��{?mmbG'ǩ��	I���	p���3�=���t�?�F�rm�"*[��±� o��V#:�/�o���e�2�R ��9�ZZ0�M��n��uh�H�p�)��R(����w����G]-L�����=���럩4Q4i6s�H����f;C�j�ߔڟ�j���!u�w�<ŁS�.# �Y���H�Q�r�I�1JJD欯���L�k��o�A:�j�{'b�Th��EK~���
����j
�p�����3�z�em�ͧ�< �7�h���!+W��E�0�Pj ������Il�K��!�ʹ3i%�}������ϟ�dd�f̓5 ��c�C���y�v��ŇuR:jj���-:=�U�����{�ay��2�\�gb������1��ib�ݨN�{��6�1ן�	���zh�I����Ho8\�8δ�����Ǐ|�7�w�VWIO{lZ�vv��W�����(-�E�w�Ԫ��m����������GK�Odo�1��}���Y����}�<����gP��o�']Æ��*��N�G+�8����Ŵk�pE�߽�t u<��P��J��l�ʓ����l�W�m��� ���������:=�p��[:�s��4Z�"B����˚��\ɋ�1���`zvww_��j����n�,B3jX�v��C����W�r����].n��YSZ���]ۋpd:���ɄV�uC�H�)��f��P�}t�GqQh��r�E�e��)��3R��Y\���'!�L��\;�|������OA�`҅��Șn��Es�CuY� tT��J���.�1����
q�(c��)�J�=��K��z�����"�#�*����G04P黧̀v��mHBRR����NN�|�	�l����U��_��_B3�C��fx�T'F���}r�u�#P'/B�9��u8"@$��ϟ[���yI|d�'��=�~���}�9��'U*�	���p���49��{¿A�R�?H�Q4�V.[k�z�spr�����?c�!�@����04��7�r����I/әw�JD=�����*�T��=��sCAoY��4{����HEЦ�?�;�t�b�_-�T���k���JG+_�'N.lo��ї���V��
{g�IRv�67cK�8MH�Gգ�A@��Z�5�/��#�'�[B6%�����,�����p���6\#
��j��t���]�(��v�V�Q D��<ڜR�K�B��[�Y�:����H�FFF�ps*�{���ў��_5��w�^?� <,c!�m������	q��RH������ȠҜ�J�}^X�0)�1���6 0���w��Up|0S�7v��;�zP�� �d������{ �w0=[�)�[���C�H��ɚ��Y�W�0���:+�(�縹��|�~ݝ��K�����f x2X�Ł��وp���*k����C:��h�א��巴P\���g�G��U<���AE\������ �q0�����5]8ڞ�m��ta*2Vߪf̛y�d��$��ɓ�#�1��Vm���L�" �`?)�6�U�:8O��XDb� !���%pi��C�����>�G2���cpİ|t�D�,W��{t�y����ͮ���TVN�����f�G�=��L�l���DxL��a^M���(E6�G�~�|R�L`Av`��ۘmq�>T�<%ς�#j�G<v2����q���vs�c3��@#w��~�&�u)X�,[�Y^���v3��;󟒝���.��|�l�QӁ��"*�i �v��O�	���R���Y^�
}��ݯ�0�jK�2����fn<Pe�WIZ���o�:��â��Rߎf��q���5% �����2�.�R���
:h���P{�wUm��, �^˶|�c3�y�$?!����Z:=�4��_��3F�Lt��3���D��7Q����2������ȓ��Ww��2Ao��O�%\m9�,�@�ˮ��~_�p`���$��n��5bY]%���~�"��_n�v��%�'0���/����8������0�ĝ��hN��w��/���,EE���˵K��L �1�*TqQS�ϯk���{Ƞ�i6bIr��1"�qCqZ,s���FWu�{:e�����P�۶�	�Mf���i���^o��Ң�.���`ԅ<7v��$%�y�p��ѻp}52�]K! jp�c� +9t=G�	Pr@����Xkq�/�wcn�:�|=vb|�Z>��8\U,):���s��)&��YJ).3�QE,�<���V��б}pb��ML�+*����gx����@��)�5��R�������h=qyjyw�X�E1��.�����w�%�p�E�԰���f�.�B��Ӥ�ؕ��E���X�Z˩�4����EV�sAx�lm���КWGp�̔�LA�"����Y�^�*2�뙼�)������ @%�E�K�V���4�}ZY��*Y�C��ذ䍞��b�K�1���r�&N��A��lx)R!���J��4�����E�?*��ʟ�����5`lR��~�	�:���*#L�D].6��l7�W�J�|�+���?���]�n���G��J�8 �����b�wm�ci��軀m����>��0o��Fn�NG��5.n\�(�}�l늄R�m���>���s��7���k��Wj?"��m��hh�֜M~��b�i���1����p�\�L�Q������^7'z**+��>�9���Z�l��ffܻ�%��$ԉبJ�O��)�qk�
��@eK�\�;Ǫ˸ij=P!�2VI�����eK�C$���'����&�?�V��:�S��t�s��U��>&�8���j�;F8̅�S��Xa��S��~��\�|��R`�������;.�c,�˵'�/�N�R�<[�������_����\�6�#�t&��܄ �r%��\a��661a��
p\�_e��z)�/�3O�	��/�-��x~_$PGc��#ȜaWG�EF�2��y&ZS����=�y'm��]o�ݫ��L�~bĸ�8x�϶���c���חv_�z��/4!�R��{7NO���~�*���:R�2j�G�����nV2���E��F1�u���#G��D����ja�0���B�.�7���8��b�y�:��P����Eo��Ea���)����h�SL\p: Ėy�R���������<ZL�t��-��YM��c�� ���}X�8m������y�k��v2-a�F8n�@�#���"����O��9�Pۮ$v����#lԮ���Ok�-~����u�n���@����"�,��%���aS�g�˜���x��I��72+Kc�Z���3O�9J��B�M�B}��M��ǌT��NڇF7��j�6r�sM��F��¹�{�7˖���F��p_���X�U�)z ���I���Z[$j�.q��TU��o�_��f�z����@]?=T���;�C�W�&5������"V!���H2W�i��d %u>�� �vp���-~�:�E>�Hߎ�X��ry�����{fR����~�|��ii:^�]�덭 ����QGF��'I��W歭|�LZ��ά���$<���
RXXȡ��][�=̛����� *�,[iB����i&gbBs����}��ԙ����xɶ�rT�XW�G�F�x=;���*��]�gt��������ϰhb�L���VW7���
@�	��J�����@��a�[Jf�O�M�Y��N�Z�mm��ҨG%͓}W�'�EEc  ��J�]ߊ��$-��~� ��?��ro6m��uUٻ���Z�8?�ցӇ+B��ڔ���>\jV�dA��n�t!O~�����������E�נ�����҈.k�w��� [n4_t!%%}&ȩ��g�8���/>���_����DRiO�3IϠ��-��|������B%��Y����5q��0��LGO���J���]�!���~?3�����6�@���S��b	F8����C�W��3U&�y���9��0o����^�x��Me�/y
:� �����|��\�-��'��VF�p"�-Y (
H��I��D���f�h�Q���$C��{]gX�"�Xez|**�Ҋ
R�(B�fG��jV����GV2-
�޺x���P�s�U�7��>�Iu�E]�{]�s�C���WŢ	G�C�h ~�E�jk���e��Y&%#���]R	���*ZY�wcO�;���pqq�L9���RCGm��Ϟ;�w����FF�u�.���0�b����QW$3*���U3Ҥc;E[]�|�`q�*���e�|�}�u�z �nS�jH��MЊ#�bv@���֬Ԓ)5t��)@����xO���n�'�[J#��t+m�n��V��0hQ�V�s�7��a�ϳsq��\mK��`�윜
&&�������%R#\N~,./aaa��\/��[q��ɉS^���zL���ޞ�����F��G=�?�J��vP�!����vv~~�A�K,��?�䎘�O�D��d�q�̖��i4�y�F���e���y�Z��lDu[J@X������ U(�{�}����p��c]��]AM���	��2om��`�����Oڡl��������[�?x����5s%)؋¹Y�	��ĿJ��p�2�K9�zS�f4>3ĝ��D��b^x�8a���0`����DBp�	�!�=����A�7&���
�2�T9����Q:�V�b�����߄>fd�Zhii!*��BBk��������N���Q�~�zX9�<�;;�� �Mw�2K������"(���BAۊ8P�c�����*`C��琛�Ln�]�,���2����a����zo�g�����F����a�\����6�8(d��۴#(67'
o�H�����/*�����[>d��I��L�j����g;ᴫ+-X����?D�\����}�<Y_���$�.R�9�:|�2���	W�V��263\X�E'��"5�a�ƸJ^M)�����f/�~�rs���o�����}�n3��e=n�"Bd�I�F�Tͪ_�w^��T������;����w��@G���������=������󠕩�8�]����^V��S�s��<������f��`��~jj�7~�į�-�LUK䂢D�w��u����S�W����Pt�l�`Ǌ������d��jj2��y�y��K�����P�uՒ�KX���b�꧂f��W5����Ol�����A:��0wR:�m�J�� ʋe-&`o�:����P酨=�ǌ�LjQqM�_���E��%����u$��Mg�o{z��/_�n�H�
OOϝ�Z��dkBe;n����yX��3�3����䔸����F���]�yo���6�1N���/I,,Gv� �u��E�B~Gyxyl	sr�iHۂgd��W������9�`��OD 0�"��7,b9*��Uw!�ĵ���O��v0��۲���Ţ6��$�׫?���q���W}�	q�JK]�����66Lt����{K>:�������Wv���Ʉ�~�/��L�xr���-|���fk�{����ݙ������ٶL/�I���P�D��.��ۤw��Z�WV*�h��T���F����~ɛ=�,0(�^}�O#�:�K��ܢ���#��Mlne����AN��L+L� ��f��*�|��(��z��f�K2�q�&⶿�zb���1�Oi�O�����na�X��a�����.01���Z���+������qH
����kxz�F),�R�t���_11}��*?�U���5�E�V���p�Et�()��:�~sR��H�
���p�O��JR�)�w@��&���B<��/���4�[�s	�r�n%s�T��m�ϮA�o�t�a^�,N���pj�J��{������|E�X� ����_/m�g�Y��%�$ڳT>��	18�����	�.lrIBHg��9} �6i��m`�R�`̇���Nz�J8h�Ս^i@�OX�	������" �b�K�ן2s�x�Y� �H�8\�����Q�����E0���������И���"��6��[��e�{|R,��v��д3� ����ϕW�e7�lX;e*��C�?��x�:���j�3�fY�O
��>5O�H�H�^ߌe����N|]ĪW�>yy��o�bi�.��O@ C�����O�$�M�8
��_��/�`�D�b������{�٦��6�JxP��n�j�c�z|��ܓd6 LǣPA�Sio���A�Ԃ�z��]\\؟�tk���5���c�{ҷ���*QL�����94I�/xJ._O1�N��D��`�G]B4�ׂ��!��92fW\25=���#�w��ӓ���\�b��^>^55{�M�::#�8h '��Ҥ��F�-�)����lt\�N�9ꤸ�ð�>�w$/�����˛{���i���KI�E���D%��Mn,��ze�q�r�O~�����Gv�@�4J-Ga0�`�	I Y�V�F�a�/(-}��M�Zo�W������RL��u ��+�������p�F����攕�����g��c��(�aQ
T�t�����j�V.l�le��u1"	�6Y��#�����䶵���I"�{��VĐ���U�j
�#��>+�?�w�9;F� �m�ןQ�"a��Ϥ�]K�Az�=�[���44S�8�fu|��fC+�w�G[��!\�#�C�Uy�?��H>^���~9��Gd��A(0��Ѹ�x^�'��O���MǜM�?��:�����+[�����0`KyλƖ�$5lW׽y��QH�I���<���;����AΨ�
Ccc}KKKe����DDu���IT�C[} ����M������-��G��y��7�/F*4	O��m^\�K��-+=��P��uȮ	5+b����y��Z�xj0+ƫz"�?�[k�@�l:$7��u|��գ����zv�Xa��B�s� >��=!{������4n'fG�r�'����bo�&���m�-0Lz:f��HC=����b�Y�g�ֆpNw,������D�5*���X��J�ҏd=ģ�mF��曟@N���~=�c	�����3r��5^aT��B��jD�������2�����w4�
�<#"G����V!��.*�B|P��r��o3��9)ji�n��m�m����,�p�#�o���*����M[WJaxe|�Lwm�m���R�P�S����?�n���ob?ܺ?�%�ϝj���~*).�I��X@.�f��38�/Y0�ҟ��@\�_�g��Q2L3�4��0���f"�g�%<�z�D�����g�{��χE:,�&��� �ujN�W�2a�Z�n������U��᱕().#�����|�������Y�.G�]�ӧ��C�޸��@�����HىW�^ii)�pƤ�m>@{��}M�ou)[Tv�	�3��B�}�� S�H�JܠS�c�$Ǫzy�!���������ē��`wlI�����3^Ա���w�C�ڏS��=��$[)��
f?��P��"v��8�����S�����<n�G������Λ�����l�s9ͫ�]��K�%A瀁E�ͦu�l�Ζ
���ף~�em�p�k��]��7D����.��>��l>�d��(|U�(g�,����B��K]P��rĿ��^rԯV�3� ݨr�V�]§2��7����׷�k�uV�c$b]^:��=.�YeQ�+;��~p@��a����+��$3�9! �����f�?XA���8`b��W]]h?ɨi>�5#~AA�b+X�>�G��^٭\�Q�43�S݅eՇB;#�i/��ϛ<6T�(�W8�q	4�e,�3�Ϸ*���}R6���H��iuq��w$"�8�!��y���� E��澡=3���:ߠL�Ђ�s��%������ث�2�d��g�,G��[����������	~�բV��L�����.D0�
�VP[+����2h����=B�Z�HX�/,�� �ܗ^����\���� !)�:����[��ak$V�cXO�jR�.�1�^�埔�:����<����3��zq9�?ëH>��*`E�#g�6`�a�.1�֑ͱ%�6w!!��-��r�X���'?)��/��������D��C��ˍ�5F.�n�ʪ�,����)�l�t�@sq9���)
�i���G�H�F�%�z']��?��^	�(�{��u�9!��HĜ{m�4�o:��d'����m�������*��qOļ%��(���Ǻ�	�� )ʌ�����lqe��]��3"S8�H�_a+��A��\��+�V�TQ�ퟩ!�4��r_���!-�J�0�G\��=q�0�r�[�iC��Ǭ,&��ۭP�l.�r��s!%S-�M�395��>��9T��$�4]~�0�@5ꭣ�ز����<i����u�'-��d\�Hxy�į-I��N�\�"��Km}�/ )z���/j�3SI�=��9+Z�i:����*V�"�[_FD�-�o���_�%X���I0.�$�X���$ߛq�R��`�U�RW��vH'����l��O
i6�~<�0K����C5Dz��_�nE�})�"�= HXnX-_��TUWW��mT�Cu�����|d>i���E�	�γ�`Ù�1)�^��ջ��p�y�n+�e�A\���ka��@ o����d.Oӡ����r��5)Z�͡T�4wBf��рR���(�_��J3�i�߇$�0NN�Z��sh�IےT�q3It���o�]�SuG���
{*P�$q�`bt4��OQ���#�3���!?o����bc'��Up�v�l����iu������h㇕���-
��og?o}�L^�P�t�Ba��B�m}�{���0��ü<1�hPZ����@]|�>7���g�������V�`(9)q}h�ihT�A��!b;V�¸�����z�{��0Q���E��G�o�^�j嗒g����T� ?����h�ѷ�T);J�&�-�4�(_�Q�Np�ny&$#��qjE:�pj��ƒ<���m���}��ϓr����.�77O�MLqE�k]�x��l��}"ږ�&����ZC�d�$X�����&�����˧'�� ^�&�oG"6ҬK�8T�h�W���
8mt��2P�E:�	��0Ul>�ËKmS�W�5����Oؒ
��iKtʘQ�����Kp��L5B%�J9wm]]�.����6�D0-,��yF�HB\E�L��p�V�'ܸ��lL%��I�(�l��dg���Q��A�A����0).V�R�á��� h�6��1�?=�QhT3%,[h{�?LPP0_�lry��u���3C�Y���d�ЗgP�"f�w���I�N����V�����	l Q\�m /ZX�]�3�ɂFT�U����v2��D��-T �����(q�6���v.��qQ��戸�!'d'��JFc��`��*t}r�b���Y! WFZ���d�7���'��;99����A�} )�̞;�����||W�b|�M�I{*z�!oG�{*,Z	M q����L� M��3��n�͟an�S��:��Z�d�3��^.���4Z�Ir�U���e�����9<�,��M!�R"����t��k�bhC0��4�8}Йqj$�U��kEJ�U�o`��I�P�	B�1ߒh�K�V���g�����ub����/2��}]��#'D�RA􈣉!�bA��\���Eh�lD,��s1zz�H�J9Ws���\�V��;uZ(j�&C#Mݞ�u�"�N{)����]��pall�_t�Rr��|0�-q���n�2�l��O���o�7q9��đ�I����a���Jp��0l;7�EƮ|�|z�.P(c!/�&��J=@���'��Ւi�՟ ���(fŧ�`�vp`���|]��V09Rt~Rt;#�BN��_��'We�`�X��pt T1pk���W�*�暌�d�Qr
�wmo�r�v)�d'���F��$�R ��nD���]**�����%g&^^"�h���"�?�OR�v�zɗO�9��m��0%o4#�@D��p��]!1��)��M��@e6;��'�`���@ӻu������w��v���`[�d�e��<"�[Q���R���<^wq�9E39�Ż�!��o�?D`�h�
�ȩ��&�r�)�Y��\@������!�IM�Z�]� �b0�bi�u �gN��EY�=����֮�H<Jr?Ԓ���)��A �Z�v�C䏳�_ogG�>G��?��`�2�;�ԽL���/�
GDv2�}\�4��(N�� ��Ē4k�o�G�����{I9��{i��0b��	�VV�WT��c3�\��JR�ddd��dWfq~=�Kb��~:~e�j��8)�
[9$䒿��+���������z4��KIKK��*|yY��ZU��[������PQ[�_�������T��¢Q�ҿ�����#	 wy��*��~w}�is�fg�ȓ��3�T����pJX�Zʼ��޲���%���fC�#B#23�|{��_�m�c)B���i�sQ����-��C6�O(����Qj�
�>��nS���;Q������P<�k��%�"K� �?��,����'u���/J��@W3Q)1�I�eA%Y���������>��R�����?��KE���Q��H��25��ŵ���	�U��Ń�k�������N��.t��L/�o�+��[�ҭ�r�����C"?��pT� >�2�~�ӊg��\��CڈW���\l����λ+N`�[[(�a�e�!Ǔ��J���h(�Zg`�+��{�b����KϬ����H7y���{��4�h�>���\��=����r�<	��]b}>�ᱣP��VWWx���LD�q�+�����_�k`q��׵���xz�ǭR��v��R���;E����/�2B�r��W�)CZ1Z��أP�m'W4�nd�OÅ�p��=�:1�P��2{X��_���.�}H��qO��eWF Sz7%y���-�.�R��.�	��'�&u˸�[�n�ʵh~����>���8im��>��Xf� �g4�6R̵��3��?� n������1#��5��i��/�$�����
=A�:F~��;J��W���d���]2�EE��rNfr�T`�\B*��^8D�75������ 8�ӳf3��^Ƃ2�ӰY��%'&�W���E�~|x���:6�eh����,������+l�F-�����5��C��ѯ?���{{{S����+ 5g8P�.��i��{O�Ƃ�C�s�Y6�Y��u�{�4�z�sW���LNY��t>�h]�%I@6�8Z�Q��YY���&&���붜�co�����?�|�D=���G..�Y�c���6���a�����l}�t��DL���ࣃe������һ�6�s.4� M��#	ػ�jc��=�r#'��6����K��H7Ĩ��?E�'ߓ��1��4F����a7�.+c!� �I���U���̉����<�:h~�X�}/��>�N]ĺ�J�����o�8�R`���G�uu�@r%D�(���f1����r+���?꼺���bK&�i�&��E�*'1�⫡����`]�n��D
�y��wRD1߼Y���ޖ�������Է[k�-t�z���#�^:a\a�HL�9_��n����c��&�Φm~ˮ�ez��y��oɎj��l2Pt����xȩ�P\s����I��n�C� $@�l���_S�7�����/���y13MZ逨��l �4y���O��h8(9+�
�w�;Xtpq�il��f ����#�vp���?N-�v4����]�l�Ҫ����I��6y |TM�d-�UX�G������DЈ�����t�o�qdo�W�� �(!R�O\) ��Ү}�����(Ճs(��?��M��?����/).��9���Ү������3p� ^����K��;-)�s��~N���(y�l��x�M�\�<�ںi�OCbbl쥢�8�ߋ�ܺ�#JX��`�����~�7uvGۄ�.Q �0��-�Fd�>�F�
 1���}øX�aS[��p�>�R���ZE[[�"�ȝ����GC,�����mӾ�[ء8�l�.0vuن~*HpOj�Ǐ�<<ۗ��  j�up���^)�� ���LL�[[Fȵ4� [W|ƙy�����m�	L��d���H�~��p�{�6�<���<�q��N����!�Ux{ַuj�yD�?D#��y�Xy��y��v
�qOm*�L��k���CK�i�8�GoNDm�g�g�sq�{1�ӷg��N�"��`�'MP nLY�J_�1�u\�h5�a���766��.���rÖP��T���;�=M9�cri�{��J�=�����]�axW���+0��{�R��G����'���4&ױ��#�|�1�xH$��nnn���Wa�A(��\�A��gm��ç�ͬL�"՝R$'+�<�`E�d[��6�����凷R��Yˇ(e�<^G�Ϋk}ڐ{�@��G�4�C�aJ�r\�I?ps�@���e��xJ�l=�X�"J�X<� �?�^���'I0[eֻ���Q�QSJՔ��D%E'�o ^� �'Ң��ƕ�_�{,�V�7
����W�s�J�U.�앰#�C�O]�)�ʙ���\��ݒ�fq`�ʁ0��'o��/'.{z0����ڵ�ǚ){��i`�. �gǕ�>E�;�Wj|k	�T��}��o�%le����<!���~����O&`��˲��WW0���>}� ��A���?D��>�O	����鞯g��� @��_�T��簨��V"H�b�V���5��bV�tT�׿�mo�����[ݛ\�ð�� ��R��J�w�M/Op���������M���g�w���T���-��pcz��҂�v���Ֆns>�ҷ{t4�xD6��%x{d7Z\��7�C�T�2~P�ݜ�O�1����r�x�y���m�. �82��c�$*y����h~.m���`�����h��R�u$��#��Qn�Hn�+�^�K/���2h� ������ݺt���F'b�=��_϶Ossʊs�Ö�Mj�&��~s>n��u����g�<��Xɖ�3��:��4)œ��l 6���ɗO}s�Mw�E���0|��ꂵ#�n���:��;�	z5�@2��-�;��ǘ�P+��<!A}�B�7%�;�;�����= {{ӛ&�)$��,@Hٸ�
ǯ�%}�w-����v�u9;Q����>���^�.�����6�p��7۶���v�� �kH��X����Y{[��#���A[Dwٰj�q=�����V˸�2D)� V�xy�-*��$ol)h����T[L�tc�D��?�ç:���dec��o���A�8Lh8���FX��A�r�mp�D,���0���&.�,�T������s}As.!��T����9�ïe?J�T1�^�Zl��o�J�e7���T��}d��Y���~����wְ��,�%8�`����;1�u���p��E��f�CVDnb|�j�K쵱����y(�+g��^q�}vOQ�.Ơ����8��j��S(.n��IB����	~*tIвR�����?o��% J�`_R��a�m��i��U)�\��� �S_$�Z��o#��B�
Bd�#�֥7y�D�X���bc��$��BP�v�"&��B�T���v�x�^�܃�h���*0GmU�U�`�M�-�`&W������C�?����򏰼����U�E��|�F1!��j�Ve������6j$�r�!虠Vٿ�HS�),,��k]�ĝ.��nM.\3&-�D�z�@}:�%� �����v�	;;V��y6�c)�F���(�n����{�" X�kI���._��|����][:���'�Jj�r2ˈ��I�����o�w.��B�$8w;J��b�/�y>�Ą��OV"xێ���v:�'.�r[�{ѯXG'��}r��p��'c�=���HGuJ_��j�Ge��	��]I�H�'�_���S��$�82Wҧ ʌ���0M����Γ>|�7s�x�Xc�&�_�����3�����T��G��d�b���<c�#����r��i����!�r�C��*j�瘛��w،Ha�h�`}b~���(�ő1W,�o�ۮVԓt �ga��<�ywZcw��gi4ڝFԕ�vy����5v��0 h���%%4?q!ȃ�6��5����g���A��o�<kk��		Y����?7��o�ܶ��m���~Σ6����q�Ϋw�	d��Tͦ�����YA�h]�����XW�$++�lo����_��Wx�(z�����'�톦��V�E����i��6�Z��lIeHd��	�R�QpH��_���T���f��cX���Ql��f�Yx�e���2l��=��5�񈬅�7A(� )���%�Us6��w�JR�7������>y��3��5�Aj��,����?�����#���������\���Fx��cڽ���iA��lYUx��|v�Uq0��)�9�KXY��K�xr�}}�J�ȩT�)�5��,�n�j�O�ا��n���5�����l�_ॊ���Z�/Ku@�f@L�J�e����n6��Y�)����M�]y�s;:9N./�.nk::��9VW��&����"��@�q��/RN�)�³]U�m�,�_G;sa҈zo�I�ӝ�O&�:4t�D�j%O���O6ېGԕ�����x��A+�{�#��F��c��1��D��N�������<�2WE���!L+
����7��5�����_��*旖~(���������}_{R��%N?X��v76�*WH��~�Ƿ�-�Ţi�!j�:��ٷ�(�B:>���;S�zB@�����bqd�5"�rqI������v2@�̿
��`�`σ`�<h��5u�N/
�����{��N4���>P}+��o��F�
����ĉ�>�z����ݡ������~�đ�&$�Az�����{�ue)�=�����.i$^AƩ��l���Y7=�]8�ۺV% �J�X6���+b�v�?w��^��w&��
NA�)�U�����ps�?K��dא�ZF����2�óA�f<?���{l�2ak2`���H0\�B�I��Iʐ�ː�F�H�г "�O����\"2�}t�җ�x��oC���B�Ł��(�v�
Cĩ���ބla,J���-�ӗ�M���*���s�9�?`I�*22�1_F�����ߓd~YYݧ�jy �lk��34d����ļ�п��r}���)��|�n��2��!��]�4\�� �Ŗć
����Lr 	����ڪ)оpr1s̡��x�Ҥ����	��3��?\�=���0��ٜW/32�>��-DE�]����$q��j�My^ii=Yrvƿ>?��b�rn]6�E'*��>n��+p ���!3���W���ĵ�YP�w�H�����r����4����w�E�	��������4��3��ţ��l�Ny-�f��kB��G�FF�=��H<_\\0���7A)���ǭQ���ې���js�gz5���7=�}K:�4���ȣx�z��/����>�H��{D�Ib��~I���@�5��_���	�^���E�������|h(= ��)Ƃ/������y�.�U�]92^���K+�2���a6�����<�Tq���0�#�ߝ������C���� �a-�	˓�9?'\霝�ҭA$v����|�yO��+�R@�U�Q���C�P���i/�Q�;�՛3Ԓ#�7M�����/��� r�Ŏ���d�Ѫ�q<VlM�cؖ'��l�Y�����0%��]V�Z3�;�>4��*|Gubh�e@ 51Lyp �c.������̶g�#���_u�	d�yIX��(�����
�5��F ��
�忮��l)ƞ72R�<4�}��CD��3*����\WW�o+����c��K�n�@� 2�^߀ ���,���.�h�*ˊ���!���0ɝ�#&��6V�S���:�v�̲F�|�m���1��!�)WB�]���˦KE�m�=1��.�_N����������j�1&f��PD�L6�	_w��n?��.:?�������*R
V�PR>����K# X���D�!m�@�Iq~u�
E��A�EzI�s�}=���6��N�$���.m�k.^��OȜ�X���Q���h���s���T2���5��g�d�{���X�"Ί����Ӭ�5X���:܎�M;<��H�*��}9�n���ֺ��4�c5�:q��)҉5�=PRw�� C��ݟ�b�R�ʙw�K�#   �׏ݏ�� h�j�誟���������%����'҈�Tł�����|�D�eI�:ר�[
ZB�	�I8<bj�x6�r�!k�G��A��lfwև�vtz�/�ʩw�� �����	iwo���g��L���`L���g_	�6t�3�~=���K�vqX&y}k�H ָm��g��"��A`�xn���� n)�YPO�曄ȸ��jgŗ�w�x��'��ߧ���0.}Q>UPQ�Q��+�c���é�/핹��:e�rz"�_D-}|��h���uj�Os����?x�~��{p�t&0,$�y}� e+eT�,��yl�%S�L���sQ)U�\Q�c������E���pt�Q��ax���҆�ofp�&�K,''N �@��tP��M
��6��=D��vIg:��_- Vc 9����h�p =yb�n��wz�_�*Z}Ƀ�����:,��yT@IQ���K�KD�Q	i\r��e	�w���e���=���{]/�p�g����=��=��[�����]
�1�&ܵ�rkFzz��f�3��`@%���Oy\]�����2�Pԥ�Y��6��KM5 l�N6�B���g�6�?������{-p޼T]s�-�}�q	�p�D)�a��^�����H�=�8Ő�J��_0N�8��um��!��� d�^y(���j�7�!���μ
���P17���s�%߇Je{�������!-S�4��Y�P`�<��xm&*kP�LX�-WcH8#4� ��oڡ���Q��La�A
��qI�[��.rg����e���r,����ޭ&�+�O��(���uH�!�;w댖��p��, ��4��|�L�����]xbbb��Ls���#	����s�'����=�u�7,h������_���v���()j-���GXkuI"�����q�3h�U9��^d�=?��JQ� ���z���gU�>y^sZ�}&��yɥS2]�m��������d�}X�[ 1��
��q?Sj�*Izw�m���]�(�Q�O�/(B_K��ތ���6SIv���<���5�qF���U��`RW7���w��U}����P� ��M��o�������KH��eΉY_jk7�;??�{�cɲ��� `��I��ష�IB�e�1��Ψۚ���&��Qy�r����D�e��prf�7���}�SSSu~�j��+�Ħ�B�
X-���4��ȭ�����gɖ���)�{K1���Ϡ�fԍ���ِ�8	�O��ا�?>/0�ܘ�P�~�=H�̠}��i4�J6�zT���z�o���6_Ru^���n2uuu�p�-��2�W���SJ��J̍j�V�&V�n4*zL�aCN��SruU����a?V�I"f@�����B��j}�֤�j�1V�nւKb�V��_��v2ݗ	.��ȩX���%���g^G�F������ߪ���n�Ė�vv�W2FȻ`˾s?�ͿL��?C��C��<d�0Tmbɉ��YȤͣ3]c���L"��B�f�</EH�G9���c�c]��h��+�$��vh�H�S"�����HY���tT�7�ac<A�G�p�CxQ�U9 �MI����Hm�c|�����'j�T)���N�L��� 4(`���R�՜��6P�X�
��e_?��	X� �ϥQ݋Z�����o*�}2�JUb�܍�� Vbrr�].#-m+G�K1tA
�6�T��a4lTr�M˕�j��/�Y�l2�*[Z����R,��շ%kH�Y����f����q�75N���|�"�M��nq��}�9��~�N�����%��Y��뱘�v� �`RTI��iE|�UB��m`��R�u ��U8�Zq=��O6�% ��N}ҖᰁI}�
����<��)H�7�ӱ��̆�o�,#�~x�z\^NTy��!`k��w��;v��z-������2`� I��Ix\��ps�$�dD��"�K��0D��������K%t�6T�߮�'����:-7��j"�.//�O��䬌��$�D�C ����N� E���׭1	�؅�;Q�C�0sb�������2��E���RQ:��;�P�������9�6�c���ɥ�	�-^�	���uy���Z-|�4�P��[�
�7[�5y՚����>N�����]��"Q���}���Hg��|8�����b|��f0E���	}Y��ʱW�:�"����QW��|��PR��b�Nw@�>o�)�������[9��!{UfY)!�G��w�k�q1��kP���z��Ub�\�XZZ^��"����x:"���(�����Q�d 2���c5K��y��s���,ZṾDj��嫉n�]"x�Oǔ#��-+x�҃�e͜�j�$0�%������rm!*�V�ؚ� �D�af>?e[�הS�n�nw�S	��������k��ė�8w	�<a"G�
d��{�Q�����ꕀ|܂���vyyoB��Fp+w;��Z��*h�Չ	�ѡ�S�%_ң�[��r�����5�h&��w��UU�����q}�vt$�O�N��'�в�KPZL�y�$�bѾxpw~J\�faJ������9�l����|��?nn�~��A�k�� �� ���LߖR�hp�ޣG=��y�`\�|uIѺ��t�
	G �f�b�6N0f*��oڔ1��}6(7I��ļJ:F+�&�/�����OTɔ�8w#�[�$�C %)��\n��7�(�r��YY=1?q=�'peS�ٸ��� Zɩ��@}��zG��:fy��J����`c/~��t�o߿�!�^ʒƴ�����r�	*�k�{tǡ����u����qhX�b�?p{H�	a�|��_'[F	?��V4ץ�������qj�A࿩E��7���G��W�*�+)w
?�0�X$��U\�/F~�\���v|\��璍�dd� B�v�� 9b�үφ�!%D4�����I�����.%S�#///ύ���U8bck`�J��@��&�dhT�;�JK�Y�'���w��g�����ꩣU��gq���Ě�g<��[_q����	ʮ	꘩��'FJl^�/Ru��泷�@Q��Zyuu����d-����%6�{�����f�qv��r7��o7��ԏaphh`&�ƃ�Kߺͮ��_������N���ң%*�f1���!
���!]��.gy���an mUBʿ�	f�s.�8�g4�����
޼�Q�#k:��PWO/�0N��Xk���p>d�>�0<x�u����0|�D�"��A����8�A�E"��4\W@
���*ͻ����މ�d)6��:9ᱮ ���������Nҩx��gu���m�P�f���=�k�WJ%� �lQ������7&"SS;�x���S�sS�Og	��u��UtQ��oE�߾���V9�<|,�e��Y{(����A�}�F��5ۋb.
����{����\��҂��I7뙼��u��V84�c1C����H��t�'�v_2�[]��H�\�dm F%g�����&u��끵�y�&��+»�����(�OQ=�����DB2���AD�����B.su|�=�g��6Hp~�M��P����P0��@��}�x�����G(X5t�^��s��?rb��"��}�yD�Ij���=�se�ɒX�V�����A�U��� �Q?1!!��=S�^>'!.7N�s��ׁ�=���
Q�60>���S]W��=�͛�렕O0���g��1�1���L7�IΕ21�4݅V�K�T|��`M�um�Sq�5���y�AZQ���Z���d~<�/zP(���?�q$a@V�㱒+�ӿM�ȏʻ��%"~��~������E�4[;����d�O�a�4��'���Qb�F<�Dߘ��QS�s���#p.�R&�2�!������LX�$�dc���2��[i[��x�Y�_v�����M�^�B˰

�G9RqiC��
ps)A��?�5��9�����U�^1��*!##2H�!(k;0����,�oh5
��ڧ+��;m�Q�΋
u�[q޽�m�n �Z��v��T�?>�C��4�oM��'Y��( �ؼ��~K�T>���H�����T�e⽘aJ��� F�+�Z�KP�[�y������27x�ԗQ�,8S���cڗt���O(��v\�*E,�� ,���?�@�:�]`c�_B ��=�:z@�'''��m����u���y�	�_��ѱ1�X����M�tN�'�!'<�c�M;~�U4T%����������t����\�`<����6�1ͧ���q��eK,`�q���f�����5�v����?w�m�Ds23���+B="�=������Q�����L,;;�cbI�`�e�\�%eb�'ͫ�E�۷o_�J��l�0���E�ܢ"�u�16�A�(���˺��#%,x��gt��Ef<_T'y�u�o�-5aŪ�_r�(�����ё]}�����}��&�r�Ex���z`8�&�Oj7���^Z��z%٥0[WG����{�HD��l@�b��R�����:�r�65y�'����)o���)�$����V���qE�D�n�<�g��|Ԟ�\7W��^<��Bs�|dW�V^�����y&L����I���ϞM����3zv�'�1���CQ��6����c���p�	x��I���죗ӛ�$�W+�}A�^���gA`|U���}e�k��)���\�W���__Q�C;��o4�+pe��^<����K1��l>�Yʦ}ZK�|�I����/�ϞgxM�Qh��D��}~���(rǥ�W^�J��!$S�����=�x�B���~��	�2�S�#�3ވr��q�W�v���[��Qj{��H�U�J5(j�C����D�{�Y�tp���(�Ec��/ك@�{gO�/}A�K���`t��8cb��_����2��5��p� �)k>���H�F?��d�Cc�E@؞��î�q��M���T,p���|IQ�)������E�������ؑ��ǫ$���cވ��S'{�Xl"xS4��v�+�X詆~�!K\=�suy�����t�̠��iG��Zlh"K `��<9�+t_���a��%�)))=�_�/vi��ʸ�����ӆ:h���Un�wӊ�deY^Ӊ�;�H^Ѡ�f:Z������S~���I%��3�����N���4�z�lv��.Y�Y����$�I�����y��|
���i�������]����:�ܟ�d�*!{Rއ_ M�|l�WcH�������Xfo�w~�����W��!�h�nd���ԾwuuE�&��*�������V7�T\�33ɉ�K����`�!k��j��FH�oa��>>��\��p_}���nW �>�*�����5SX8��&ߤ�}gOr��m��
�x���-��}}xQ ���^��|Jg�"�s� <���Q��]�-��q�ZJ;d�cƋ��k���"a�Ύ˭��+����1�����w���	�̱�3hbrJ�?:�\�g�<w�%���TM�Sm��|���4i! TW+�i�������jf��@��E�.o�k�G���zؽ���F�e>�,���K�I��UB)H����1,���u ��iO>؝kkGtA������zҀu�1��B��h��M��[r��
�,��������l�p_��
!M�3 r��������Ն��U�/��%�(t������A%9������m��c_����C���P8S��Tml��=Ne7������Ի��M��P�	�����w�Bi%ʩ��j����F�g��CX�q3Ed��TG�-�d��}� �m�!��a� Kַek��������e]�p =1�\Qm�W8t�N���<�JM��.D�a��Ƚ�i��η��M!�525oa]�䘹�O��c`Y���X8���}NOu�u��p�G ���XUM>\\��4	���L��p1` xum�5�����OF��7ـr�w>��)Q�F1�ȁ��yj�K���e���JMs������+�P����T�5�~}�=
�˚��\��`�x�f�08D`�F�Q�GU��7!v<�?������e���2�q��%��M�򱉙Y|��C��z���m�gǄ���xٮ�к�z��4�C}�G�RIj������l6nz��H�W��������~�����{z�����%X�BBB����P{h�8bfFzx��k�4tJ���2�`�if���*cX�?�T���v��0~{azޕ[�1��/�J�2+��KQkwg�=8�no����zF�'>TǺG�w�o9�x
���88�w��1�/G$��dx��@4�0���6�K��o��g�Iz#!kg_ZT��f�2C��� ����
��hi�����&݊�	XS%�u#��4E̩�l6� `554� ����H��Z��ySf��F�I�^�~sXe��L�U0ر��:/ӬToQN|ʰX��v*$}�.��n����l�?n箱����v�����P�cs�E���O���͸�ޢ��܁WbJJ'��އ��	[�#I�G� ��jj����A�B0L�ox�c��������6�",�"3�r]����:Qk�����&a�ܒXNz:��������1���97�7`��q~:��9�1���C6�"%үp������I� /RH1����|`���Ξ%�mS�����ez@�������.����A�ڝL�����<"3�ʭ'"3���D�?O����({{KpF˾�����f�~��Ȍ�b?TWW˦��ų�2)�"���<`2d���$��U�`�l�$ϟ�S��z5�1nĞ#�I㱔�i:f
�����N!��~��d�jF�A@''d#X3���M��2�6t���ϵ��P s����ێ]U��1Ŀ��ǉ��7	)$/���w�˺��L�l'][��up�*љטI�sq
�˗��5(���Ћ��lN'�wj�7�����6�1)�'��RCS�u��9'���=��oj�[w�`��Q����#��Xx>,Qӥs��QY�W��{�Mk�G��>[�T�5��<�v�z�������O�8E��Y��Q��}ځ>��V����U?pib98 M�߁�ت}�k����=ws#y��gcS�+N(`�>���}�O��������)�<Ap��V`fq��3Ar�������7�b��cU���6,kڞ	�.�KF�,�Zq��mW?���^ޫ���R�xJ��O��+�j�WFA�T�;��������~�L��PG7�y���%#y����bfċ�Ý/N��Z�k;y���M��++V�����@��WV��D��������M�>����-���]"��&	�ŕ�S����7~�7~M����م�ݬ{IS:�ׯ���T7�ז�ӊ���s�"�iM�)%܊	O%c|�68�(\���膒�a��S� ߳#(H+@�����^�
�c6�ւ�^���l�O�h�YVMλ��|�n0�/ ��oS�c�_^%U*��:�=�-3�[����U'Z�J��ppF����(�8]8�fU�Đ�n`sP���xFƙ��8Fmk��k�c��k:������v�_w^^޹�#U)l��ފo��n! �Α��#������6�=y�tvضȜ�oe0���~y5�f��f�$�g]ɦz�1�O��14*iֿ ����s��1Vy���(��|I�f��H�.����n�p4UV�2�鋹�7u>%y9��h@k�����\��Y��͞7^<��2s��mׄ�`4�Qz�{�79/�Y�0O�e.x�`4���u�^u��\6��J�� ��'�t�ߥ�{�U<�kc�f�3�S!�P�B�z%�ơ�9�������O<�J�CC����U�23�%���M�ak$��^�O��ў9zI�Qrn~�͗��L��O����v߾Y|�����xOY�\�
���\��Ý�x�61��qZ���*��~|d5�b-%��n&��陼=�uo���Sٽ*|��ݠT���� �mmr�S�w�%�{�BG�GJ,l�Z3��?M�xt�6�*|��� �u^܄���{�jK�Xy��-�b+���`b�G��?^P�;=&�\FV����X��`�	�Xc���O���-�/H��k��5�����k$4vi�i����>����2���F
~<�gf�9LBFF����l~K�c���g���7����p��s�[0�bS`Ƈ�3�������6�͏Qƥ&Ȱ�v�����ͻ�����O)umy�h�ު�O�>��>
�{�O>i�7{8�{O�ߴ�&s���r`I)((�ۛ���F�V����+V��W��X�)8o��e������+��������l�Yru>�-�&��4N�((+���=���0�y֋��Y"�����#�yV�uy?'��e����;��G���$�ٸ�'�K�����ʽ��L�eGq:d����|��R$�l$�2�\|�Mu���Xx$�!�'&Ҥ0�!��/"L�%���8�j�?�w/��#�ۚ�Xz��0#�uk����N��
��~�BK���� �'d�=��L)��dh�(��JB��*���ӟ*'%UB�����$�A�����6�t��;���!{�0�Q^Pl��Z����ڢ�ѝ�X��/߾E��u,l�Y� M�o�zԫ}� d�����a�h��ձ�R��lQμ1��M���EU��%�1�g6vv��AZ4��n��:�bx1�<峰��`r�u��}J{�6?oȻ���7˧M<�^�%}��e�lM!`l=�x&y�;��8Ym��BC�U��Ŭ����Z��yե1�(��i�:f����6��eo����Ѭ22���5=	�u/jo��e���,|:�����#�ڧj��bY��i��넌�;�e�l��{�jڱ���.�=��Fϔ��-ebx���UY�V���"
��v-,˒�k�P*����E+�?��G�7���-e�z��I�[[#��tI|���� ��=ǥD��CD�C[��e2�e�L�/E,}�NJꭹNR��7���̝�=���UmC�F-ރ�������K�T{98�Y9j�f�����+���2yJ��&�?22��W/3�O�I�H/��I!'Rq�;ۂ]��r�N�!O��'&�)�+=%��.HoG�uk�DOL2�E�	���Q���V��Q �\\�ר~q�L5~��߬�>��Pbx�$���	Y��݉LYBG i�⩛�z�]�����\���-Ur,�WHvI�_+��9����S��ӧG��W�rez�	٩�a݌�hޜ��^�|6��a� ��s�~��@�wƞ���ѻ֪����>KK�Oj�D��9���ˑ�;`�=��{~�^��PY��uqEY[�*vvF�͓3���ܟ�1��HII���}��\�ۀD�ȇ�1�<5�� �񄠺��ls�\]�}-+��f~���rf�=�{�:?3y�|wY���tbr8j�'�swc(�U��s��������g�x�����sꖧ���1	���1��Y^���K���wb$RNI	_���fs� �xn�(�?Fv'��qkݬ_t�T�?u� +C6��N�?ꇾ����b�W��������g�Y�0��#_��?E�8���ݔ��Ec˻��r����_��aE�������\��}�=�뭂����s��
6�E���%A�s�	r�	L��W_����lx|<c8�Y��^_�~'Xi��I�n��ؔ�1H@@���l�|���8?��,kۻd��^x�������[d��˵>�s+��"	Hår�6P���Zf��"{ �&�]�zfgr� _j��/7�`9R�T���=�*6Q�ium�;U���***�1<-�ӽ�s@m{M{��D
���+���[���6X��m-45M�[���!O!�ug�0aUERS�1;kT3~!�g��Vu��إ�3u5bbU�Vp����s?Q9���G	�5
V�l:8nz1`L\��hcr�h�oi%�Ҟ?�iy�m�t���zkG��ZNrrpj�-p!<���ת�r��:�mY�b�g�g[����iA{ﺥۆ�)�I9xa�G���$d�	�ˉ|�)��2߷oY��H���^�N�h]qG�;����0�yR�~X���v`i;I3�	��6��T��>}
_#$��Zs�+ss���yww�r��5U4J�:ښ��%7�T
b�MVL�
�����q��طoر:����Ҙ8`�ק*�=^~�˩�T�O�-�Յ��_�6��S�ko�gv����˨��R5W��T�n�G��:�.�, T��dq9����\�r�`��/�Ht(B#w\�]��jk� ̍P�� ��J��iD�2�p̃�C@
R��)��Q
�-~R��+���-5� \
�ܢ:��	r���0��yTxЏ<^��/��K0E�R���m���JԕIep4��i�d�o���J�*Gs�e<�ޯ�qY��1�H+�X)&H=9�j�����!�=!?�"�Q_���n��J�1~X����X��6U��X%֨���?+�l�j|���ubeB� -֊�S,��ܚ^��~;�q�/�So�Ʌe�o! ������[����eQ��|�mjt�؜rs{T][�+��R��H_���������s�y�G�`��`E���2@m �(����<~U���D^�E�j#�i�Y�u���?�/41!��OE�5����ߗJ:((6�U6u���N�Ĳ��cd.��b���R�H11��׼ *������N6��x�����������Lm��ϟ�[���׺�,a��L���4�E"kkȈ��~�|��x����˯��ʐ*��N������%z��N]�:��L�_�MlO<qO?�Im�Ԋ���⚚�����ʻp�0���U+C�?[��j�u��q����ב�Ҍr���];+֟��{�l_X�B9�I����`�=�.}��3:�����D�Η�\rŰ<�u�z�R~zf�""]5��j-d���y� >*cck���ɷ�֕�H:k�xc�v%�iP� ����	�ߔ��Ņ�����H}[b�`�s�lM�w�������Oɡ������e~�T��ږ�?1k��� *�ٲH)�a�n�ˈF�_N��Ř��m����N�BΠ���g��b3�lW�QK�K���r;�
:l O�-��QXv=�9��:\� �_o\��{ꗢn���?�o>i/LC��_��~v�����ɛ$�d��4�̦Bt�6c`F��c����M1kI,wJ����`C?}�-�Fe�?$������˨��}H�>� -&Xww��M4��i�0���3f�-�fW�uή�9�{�Ҹ0Zc���)7'��~uz��&�:�6���(���r��8��a��Uq]q����m�F ��.i�)%���g8dJ�6̺{;�P
0����q�ׂ��s��rrX�2�h���_�&*^(�O��e|e���rh1G~����_�u��6[⳼'�c���b�ɡ����$$yl
O,�zH΋�N���7k��� �cg����1X���V�(ʏRH41%
n�(Փ�۽��ס2��x�HaC�ґ;b3�w�����}���
����l�♽G{D�x��
^�~�#s&�C>��VsƯ{��j����.`f�Fw{q���ތ�=O|�B�&��7�s���8���6V�ٳ֭=f��Q���T��$�m,]��ư�ގ��>���:*QL�Ut�w�0=N=��l;�����#�$�s�!ͽ6W�(BO;����9>,�vo������b?|��giqn�r��u���K˘HI�	�YjsڴԆ6o�/����H9���%1���ي���D���Y�9S���O^�EV�V���J����]��`)�h7�}k1�J�&v�;G�����@:�vz���lb7���|[ttuu�,rz>`+k��c���%Q)�Oh�11̷rZ(]�@��^?7�4�`��hػK��	[��g�Amm	�w��1�K	��읯�6���]�|t�J�.0�ZM�T�8��r3��1����JU��
�T��e���-Wf �\�yd�"BC|;4�e���	И�u�kpJ�hZ�[����B-��LC��X�yA�ӂJ+ �VHd��,����B���z��~��$�g�����K���x�` �b�U�~W��ӑ��!_2S�>y�������!$v�K)��.�_V��X!&JE1�a�)�Go���}��Q��x�\����6*�������~K�Q�[2W���2�!�o��[����+>�Qp�p��F��t�X?�+�x�g��4㏧���)��;lٮQr����W��

�e�����rv���2�냃��V� 8Yr�EJ�����yo���������r�>'3�o�����9�t�$Q�{��U"�a��Wյ�#b��Ǻ�Nۚ�
��*�����?�MDEO*�7��7U؂�0�Ŷ#�$i�h��7�f5"N�\���u���2X�,�۫¢�rr��*��)y��]@�ZU���˴���,M�HN�H��1��?���s^٧=��%��!��K!�jE�{J����P��/�V��>m|�t/�q,�dU�����}���=�hE�$Q�����'���db��n�� ����A˝=kR[x0��1�W(+����E���N���ч����A�����
gS�t���4
�ֵ��:��Ҟ(%��6Q�M���j9f|�f����+k;��}�j�f9��mu�)C<G���pu���S�afL <�v���E�ۡ�R����E+�۰�_�p���MJ)�m
!�z��N����Y?��йS��T:N����vl�/��YT%����<���M�c�I���aꇖC$%J^���y�p�쾎�Tk�߃��cw.B��73���+�L��qLnA��u{g_M!(?�MHܛjA���v=m�{W�O�$t(�,��g")��v"��N�5������Q^w�>�PYFY[=��B�/��;�-_��X�e~�L'yґ�~��1���'�U�@!�('��< ,��5�4u
P*i�ޮ`Ӛ|�Y�%$�S$���y�AN�����͋���>A�q��Q�x�}<��󙅍���g/gR�������yW?�EI�q��'G<ӝS�ş��u=zomMa�A�F_�{F�C���\�X���a��.q��W�X|���J�C�{<zi��JBt�a-�ބ��~���\< ��顴�u옓��R.�Q��ȍ�z���(Җ�t��ۉ����P_�5enQ=y�ȮF�t�QmE����sIU<��S��D�zu��Fv��W��y��_�f%<6�4�f���9���9wR&��{�a;0!a��jdw'dld��ł7���(�om�kc��{}�a@���+..>W1iQ�R]c�d1^��������F�dx�*]�,q	<����?��鮛Y�_
S�D=��q35�/~����pD�DB��T�}���LSf�LLR�}���i�.w�x��V��|CX"**�B(u�ݣn��G�p���G�����X%�'�*p]��6M�����}�Y�2�ު����z�(x�~���'�sʶ���H�����J��
)��q�^�;ʖ�oL�=+��Q�<�+�#�1#.�0BV|M�-v�n����`!��px�]��&-��Y*�oA)?KB3% >M�7�o+��+J��#�	�Ǜo�jF�)����2����P���*��|C�2��`�,䧼��K��AA7$��0	��7���su��D��c�)}Y��wX�x����U������e�1��"Ֆ0��уv.̽B+���/S��0�����A�&0�e2>
֔ے �>�'�~���Џw��=��I��WL[)<Y�C��+&����"�_Oҷ/}R��:�����TUG2] ���i�Ĳ̯d3�����vB�kb����:����{��>��
.0j�2�$02�q|�;��!�����N�J����R^�V �'a|&lC5�)V�M�0���jAJ��r��;�d
{��oÅ����I �\��o�Ԯ|/j!�V#g��l��*#��G�����ޞ_F|]�?�&��"��C�:���յ�E��W�0�*o�wZJJ�X�,�t�t撷��f�K[	����_�/-���=}���iUdN31-.����Ԁ#X⥥���O޽Y�E���4��00�O_����6��V_�v�"~�O��Sx�����z�>XF�YYI ��5�:�}I�> ��P/{�}6$���CUI,��0{s�1�������t�Ѫ#M@s�W�e���
@!��RP�N���}uM�5���:��;�qqq��k��!ѯb��"s��	)%n�k���Y������M{���E��0\�o��Q-q�����_\Q�V+����]�dDU
�&���s��}F�(��`������j���1�/�)c�Xqp�߾��D?��|5������5�N��m�/��`��������#���ջ�Q��_�|\x�L���,�W/�;]�xv�)��02�����IF��r�O�}���H���}���Xި�(���J�aa����j�:C�����pA���ʹW�� ��}�W��Us�t��iF��u=3�~�����h��q4���;w��1����K�&8���3Z�+�	w�שဏ�lO:��L B�7i��#��<<�Բ��e�.'���MG��u�omlʩpx���02�ZUx�`����-���>���M���߄Ka�I��q9zԽ>#�-�W��W�)'g-��&?<
4ӄ4��27��E��P1�A�[9�;�>ױ��ţ6o������I5��K���88�h6M^����S%��;;�,!��'�Md��G��\���A�,�|�h����!m�c6��=�Y��ܮ@(u���ʪ���7Qa��o,)!"���Z7��"/>Z./b���^V�����d���]�����|��G>y)�Y�w� �o�Ǎb^i�[8 �Ѣ`&PBM-����y�>��=D�N��1i�_�:=��!�o�����'64*�o��4L������Z�mx�B e&�J�P�!��#�7
��NL$�����5�u{�|?c(='��eE��#��DL��D� :'�Ί
Pz0D		�{KK�r�]�׵�5���y��sҩI3d/K�ca�l,��v3�A����(-=e/��l���,����KM
1�����a��611���,�k�a-��&1,xTh����ŋ�YoٺuԢJ��@�n�A|ݭ����
Ș���"`�H�|��o��G�DgI ��S%�����"�kD"�7�;9	��2���8_ܺbj;Qf�)���@�c߿񄙉A������s��5���{�g�s��Hz�ѦE��8�0ݠ���v]K�j��C	��5%��7�����?�fQ�02vM�I�sЎX��x>�� >9�v��z��D~>�kPl��=��8�p&�̦��P�\����d���(=������1�?�,*\���ԱV��0%����;Td�ڨ���W�n���''Z�yA����h#���	�v&J���}�������W�TW�\�K���\$i�9������5e)� o٭y���l2sH����|ܿ-���e�eѢ����/���`]==��=}}�Դ��=���=�Qz^�'$x�e�m�����l	n�N�M��wp�{k����Ag�i����]���0jN�[�(l��R>�t9��X����W����0�v�t�S�q�
/7�g�իXR��y6=��Waii��9����"���K[��ܷ�������T]C3�\
��އx腜v�����xB�jrB�P8��픕���%���d504TK�z��b>��F�*Q&$��4�7��V�BL���w��d��,)����.'h<�A�jAl��eC��SԵ`#ԃ��ً�;��$x��}���?�����}�D�ٳ;�cA������8O�ѿ�mZ=�/�hB��3��FK��º��W�38Œ�9=��4 #[���ªV���/ GG�uDJIHɳ"���hj�۔��!�J�m�-�o��`�#��[��1~=X�o�v���D>?ś�9�czkg~Cs붾mˬ�W`����h�=bk���Y��w��,r�����W��z'�0z'학����p�	��%nh���͛76[K��2g�*�@���� �	��=Ue�]�{J��8wr�A�R�C�Ϸ5�%����&U�7gq�ʦ�������Ry�e~��1�+��#��o��^���,ً�|ی`JQ���y3F<��P-&kP12:j!M�u-'�8֭	���^���5NHH������:�ZD������wEe�Vu����ß�G�����FN��^�ȿ�
w���ϭ%oj���"��z�PC��Ou�~0�c��V-��TJ[i�2C��kg�h+'/.��-�y&�rs��ֹ���*���5U�W`Q��V~X�2aR��5����pvU�~&Wf�}�V�c͕�|��.ӭ�|5�-���Z���>�~^랤[f����9�����AT����X|���$}xJ1�w��9��.��Z��^�u��s��7�Z����*�q3>�b�����Pu��naϹd����Ř�L�`��J�H�Ն$���)��󔄥�����V|9����񌻦�rF9�� ۠b`�R83w�斢�Z,A�b�kZN����e��x�+�p�zs|�IU����D�헍�v�+67Dc��08�Z���"0+:�{j��m��^�H�LI�Ř���i�j;WoH6�(�ꧾ��C�[��j�0�D�O1A��orBt3�<���z{UqaCO�x+�5��M�Z�Ju�Z?vF!f\�2��^�����XE�c`e�%QhM�-�<�E��2*����� $�H36l��׆&B��O|`������!� �nL\�쫗�|<���p��՟�ܔ�������_�wo�2	3��6_���R`Uc�DZU
��tL����W�"�3eo���U1o�<�d��y��u�R!����?�������`z�!fm�RV�j�Q�M��"�]���σ��i<��ՍM��{ �z���~7"��~�����;��lpM��Zf@T�׫�M2M�V<T�0���r�ɷI�g���' ����/��	>y�;C����&�����;Ɇ0�"����y #![��!�Z�6b���؛h������`,��U���	� �~�P�O�T��(N�A�~ߎ�?d�&�W�;'�( ��ƚ�p|��}s�kBK-%�!ka��K��7��Ѫ��Xu��;Na�z�E�W�): d��ּ��y0D<��6T��0���'�xFz�AEaggg��%�N�Gw�`/*ԟC����z!����VS��*97��"|N�m���[�?'vm�d��A@��� J�wƮ�'J��.z�RuFe{���)	V�,��Xß���?�cD�V�0P���'':�<xx���Q�El�ç���P�AK�'�91�U�{y6���*l�$�ck��1��aQ�]�0R")�% ����)�8t��H��C������� ݒ2HI�go��y���뒙=�\k���+X��混?l���J���B5�P�0�rvv,���o�I�n}��?� w-;G���gq�c�#%e(�za��Y_�TKU�]�o��U[l�a �4S�i��������F�A�A
��F����Jt�>k��K���Ħ�(E�L�-}f�Ѐ5E�7}��se.�����]��9Vϯ	�c�6'�z�ؽ���cV��E<���V�0���x(!y��%�(�Y\MV9ƣ\��<'y{����`ft��QL�ᅄ�=-m8l�#����SN�ZZZ=n�$�c���*E#i�L���V�`�H/>7Ta��\��4�X�8�v$��:>)��[�ǳ��Yf�����.Ѷ&$�y����H�w�U�ɻ+��&�_T���=�Rġy�R#1����K��F���X�'/���nz"��<E�Z�ز6��i-��7�8�&�U@�<���9�7; /"��O�I��k^̹�{�2��~�i�7?��Sesx6ō�}�Er}��I
���2��ܣ#�Z�z�x���*�dܘ�z��(̸<;hkgc���L;��t`m~F�ִ��V
"��!����s�p�Q�eI���pWC��Ș���dv���M�<ט�Qf�a���G�����^-.�P���}x20ǣz�/��i�؃'?	�*)+���MI���f0��4*�J��$9��Vʄ}̹�v����z���x)p?N��L�Ͷ��7�|��_�Q�t�t��%v�%1q�CҼz�,M0l�$3y���K]���2hų��)�$�D�aѕ��6���+�^<�U��՛����gweee��999���[7�H"_���M�7�˷4�I ^���4B������q޿x>W�)*�	�)����'����ƿj��Xv��LQ���P���t|�n��Ȳ���#*�z�n�Rbhj����t�QXxy�¶jMB�r��;��{�f�Y�'ｽ�v��#h]Υa���-�bhno �Ӏ(���4MU�Gi���a�z��Q�B�0F�jp�,��7�L����\[�e���_,����w�M	ê��_��hS��hn��XX��s|�,�^�"Fhݝkk7�C���dQ�οؾnam�%�N�O��� �z f�����ۿimq���྄�z��Q����9���FW�( +�aQz~eZ]^U� ��$��=�����`�R6���<;)��vfhW�.�)��nW�����V���@���d=��lk����՜DG�&���'�6w(��G�q{����M���z��qܑ�}.�Zuuu±H�da�����K��j���z�9嬹\o'7u ʅ�/��-�5\���Ю4���X�!������0%m�����-�E㫿:���>z����)x�Nqׅ�բ�!*��e���6}�)W>/�v���E��.�1s�B,� ��KK�nnn���Xț�3��$��_��������0�2�����%a�=�̫�&Qڕ�`6����w(�W� --���o	��k�x���Ѳ���d.l�����Q;�ԓ�N�	v���n<AA3��r���&���0���ܨ�V��<W�{a�kz��e��h.$�J�}���*ө���������=��<�j��@�˨[�p��Y�$��8u�-Z|�鋒�S������Ʒ��bx��泔k}C�'���SiF�q{��$#���Q�%��#�\|���� 7�t��a�{��Ǥ.'�dz�IE���s����AX�͎���DVs ����Z��	Ģ������_�g�<�$�o����C�,_�]�4^h��G�.WK��=�{l��ⴅ���lԁW0�ٕ������v��x,Y�A[[��TX@�����g0c1k$`s��R�qS4��u���ֻ��@��ׯĐ	�����rw�%�J��ǧp�>�>��X4zu)Ӳ�����+(}!I���H<.���;�x�3:��g�������
����hP4���!_(��C�x>�M[�|o������9����������(X3� @q9���/��ӌ2q�r��	�%u	R0P��7Q��è�}'����,n�i�i��cr"�ۃ�����+;��ÿq�ha����P��v�k�vW��qm���`,t�B���~����ƊcFs�{/VM�fc�����|r�6{E:��n�E#D�����a���wuU���D��ɬB�W�����u�1�`���OknWE���� UƂ/��+�F]i�������\�bQR��{8Ap �����)�Zx4Oē&���y"RPPP�e~o��h�e����ohk%���>>;�0�Eth׹���.�w���N�R�,t_�	ll�@"Z瓹0���q��ۏ����^<%>��C�E��P���%�_B��yR��R���UOj�XA��J��ϙ_����dy�k�8��,�,5��R�p�wv�� ����B�Yk:q�%ytb$܉���BB6��T`B������p�<GU�A����܅���e@_����Pg�*
���r�x�4���6_��#U���>����D�j��V�����s�e:��-�X���ҧ/�DyxE�۱H�5�!��<7�}����{*⦡/�����x7o��e�?}�	a���,�vd�^�4z4��8���#jW���d,GZy˾j�iI���}��CDH8u��V��sψ�}z<#�F����>5#���2���N5���%��3�*٭a15 ~����m���`�����H�H��qxxT�?mK���Yyu��է�J
�����G|I��=�|Ż�'?���βDC��ONW�3S&�!����o��B���E�����;G�W�
��xf_̩�j:ډ������\�pd�
�L���Ш$��ǃ��2�D�;`���榆U���5��%���!�W����WD~��9��w]�A����E%VT�+Uo�����gr�vӫ�~�G�h������2������VyӶ�������u�+{�����ۻ�ES&�Z�A��_ h��Q� �a�QM�H����y}��sȣ�3����7I��QV�9���\�_�\��#�s�Y�|��u�y��V;i�z���y�w��+T�%W;>�����Ӱb���"��Wkz��lrdx~9BB����8~V�#�<�kq�&��F����Z�TT��ϸ�ct+��r���}�5}�����S����;��>:�ciq�hhi�'ӓ���������qwe�h����JI�gQ��&�f6�'Z=�9c�(�47��	ˌkFu��G�3KX����+ށ1
X������W���%��ۛ��˾��xq�h���SVmKӘ�?.���I4F5~f8)J"P('N�HHH�"��TK�Z�;��)���+g����A��2⸠��qT�\��la�ۅ�Y6��H����P?g�F�T�2����B�����]j	��,o(gaaAM��,Q�[����&$Q�zwǠ�;=������ŏ�A� �ޅ=,��iX��Ǭ���bA���/bb�h��U����X\��-����L@B00˧<%W��?�!���e���%�)��5ٔ�Op7|P�nM&��Q� ��9P�x<u6m�۞�Tt�&��m�2���1 ,��x�����R�y����ޠn���,�%=��J �}f-�F������g��3���d�r���V����ܷ�>D�`�[i�1w�?����}psq����~���/Xc��f�c�ޝQ0/�&B��QG'5h:kSSCgMM�ǜ�H��O�>���qrrj҇��5p
 �����Ƣ��di�c�@!c)��(�⵸a�Y�~��-ՖEG�����w߾)562�/,YʧT�-��p��b�;��CBL�HNN�QQ�W�z�MD@���'v�v:ޑR�o�'��Y��px�_���1�+B�1��!u�!�/:�1i��ki�;;;��������H����G O�~��}lxpd$��7�{B�`v�1]�����7c�)�fR���[ZZ�?�!��������2��E���j'�z�G ��7}�0���\��,�=�$���OID#�y�L~aa�3��{⅂�ďa��n16��w6��>0B����>��l<���dqN�ߔ��P��
��>s]ߝO�?
H�Ύ���� �&��Y5���瓈0o}�Z���j�,a�R�Ik�����!����v��ō	$ ��Cv���}��U���?����o%�G�I�.�5�3R��q��>X�N.Zmf\1�o�TN] &Ƥ@�r�o�{��	|�r�,BB��(A���|j��R��a�#�f��7�U���*�f�G�L|�'S�h��]x���,Wf���Ǧ�(5yȸl_��t��!�$-����&�0(��X{#r��*][�6����~����L���%#���"����]�`�-�I���5p$�e�yݖ��ҝw��}��� �o��yt�]ȫ�e��m� :�:˓�FI
�'$؞n��Ȏ&��8��kt+x���2�����i�}�_
��y�m([��wě�L&�aG=Ǝ�)r�Ϝ����~n�N���;�+GW
��Ou�	X	U��j��(;9 )Ӵs�ve��A�
���$E���7m]���'4a�H��c�۝��պEU/�u�#!bB�3K^�=^��c�d��O�K�9�'vo�\����������4X�L~�C�qO�';�ͅ�x[2�Ȕ��_M�����w�����:�:�O�Z�P��#;{}|�K��ڕS<T�#K��A7C�K�ibgK��/)��D�Ik|,R6�S��J�`�~�@k%k��߻����$�$S���t���8�S��&�:�:�����W�MM��j_J�ŭ����ⱆ��
@a������@���?�R�'NNN�c�f�>,y���������^]b�txqn{K-�SQ@�l�n���[�@����2����
�7S(F�{����ܓ��*��vV�s#��>�b���V���r!
�&c�P���u������;_b�iM���">������B!R�NN���λ�F�bĦmn>�����7�G۫%����I��j�g�G��:����L�#d�V���yAm���]Ĵs.«�w' ���U�����m�鼤zE��j����x<�@���������R=pb�	��!��͢z��N�d��Kt�9�Td���	%�ʵ���,cVο�q�_�;���c^�������$�J?Ω(<{q��jN���X�E�MF|ϯ�d��ĕ����\:T���qp�w�џ�w����{6���iV�?���S������j�D�2�+黓�|m���Ќ�W�Y��UR�h�fPg5�`؊���א��m(���H��\`�=�r�S�&H�1 [��Q��|������6��,%4J���e�ʃzc�4bbGWW�U��Jk�&BIĀ� t�=D��԰��Y�{%Ɋ�-�w��೮��n�m���H��[��\׻���Ou���!�"�U��`/�(R�7�Ao�}c��6���'�R�7���;ۻ59''�~Ʃ����0ү�s��4�ȝ9�A ����/���u6���\'i��Pe|\@7�i��}%g�CxԄbp8���$ �����X�p��m�(�{��b���;M�(��6���:���::�i�� �5R�!ѝ���3ҹ�b�*B�	�x0�z������D�z�g�5|>�VQB:0��U[�k ���'r/ؼ��ƴ�e���aEK��t��O4"-/��'����C�2|��6<��O$%i�G9q�ʼ����x=4ǖ��_ԙ��[��U��F�!�*I�ؗ�?.���XJ��_x�W�ܿ���W;�V���c&���qep[2��d���pR��]ZY�Ի��{�l���r�-,4GG#�c�=?�W���-r�}?���l(��J��[9�,���?�����W�k�4�1E���/82�������5y�U�~uu�f�e�&�ܓ��%EEE��Q�z(���I]��
f-'IRYC����ۺAEf$%r�_:̊�KI��s�ݰ���<���\Z]������F���1$��;N.K*�C$o�t��LK� -A��II9�����(6�_O_���;e}'�fDI �KR˭Ј`�{�*�svf���Vˠ5Ŏ�����ve%ƀ��+�4��$�v!<u��T���%�>6��Ym�Z�ڎj�
��g���ٓ��)'jZ����Q��,,�0/����L�7�
�glK�$2T��thX>�\r<�+���a_�΢ <W��LO�ͮ��,��.Vs#	U����w+�H]N���}Ζ�r��D�L��_����bt�&��4�Q�x���ٰ"9�]|5n ��#�����Z�����k�y�:c�������og{��pW!�FW] ��9�dm@8�q& �A�33���<O��\&�PKǮ.5,d�=��9��6Wŗ[5�,�u\�~QӨ�-�/Hy��sm�Y{�m0;W`KaD��(�-B�>`�T@���'��Q�9�O����k����F::�H3�ՍC�ud�p�FhτR2�+���n�\�,='�����~�m����z�����ȓ+�����}��I�Ȳ���=���}������=%]Ѓd��� ��p~~^Ui��Vo�`�=%-�iG����y���%Mol ~� q��
p�s����0�+�q<"<X�M0�=UЏ���(W��ˡ���;,^��kV�!O^��Y[Y��_,��H{m��ߞG����V=��ޡ�D3��V��K4�큞�)(�N�n7�%�C��FD��R�Y_���mQyDB"0h|�L��\��� ��{w9v�Ɨ7;�P�*I	�h�ʘe��qm��S�F��б�O�.��
����/�ha"��r�h���i��Ɛ9��0����/f\��L�i=���`)��VUk���VEKkJ����������|�ܩ�;�*[W�ʕ�hl���q�G�nS����C݇�K�ܖߚ���^_O uL���߮%����*�W���:����	�����e�v����+�Sh��5�������{�v�?��\ʄJ{��oaV�x*onN;���J/RG����7U�����ܨ���������Ǵ��b�Ր���JB�!�k���p��-�b�uC�~�;��6��󾿸�������`1�а��+����f|�vڂ�4�Õl�� M��W����v��FI �*�����2���Q%��wAݭL��-��Qz�?������H�6	n�����y3*"� 4��<ױ��,��N��PQE�=70���� �/�pLl�U�+������:�r���y��ת/�\�C���!n`�mشR�h����⏱��~I~	F��|�c�<wЕ�e���*D �I@Hpu�\���F!�I����D�h��:��#Y��))!��K#kgw(ʘ�5���q�A��`�Zw&WA}��TZ�4��<�W+y�>��G|�M��L'|w;��+%�T�n�������"�'�K'�sE^E �V���ki��s~�ʁ}�Z����]j���m�U�&�W~-I���ze��9�݀B�-g�,nT@A����!��zD�$����������je�+њ�j>���#�*��Q��/`�Ʋ��C�S���U�M��*4/��h��_u�����Ǥ.24oZB��Zh���i�I]&'�<�rD�p֢c��b7���D�p ���(���d�7D�MM�M���s�g%~���|֎�>���zV,�`�}�HI��6{zak+e_A֘>������.��s2�S(w��qxh�)-�_0����2f�Ē�@�6��%`���Wַ��|PX��ok���3
hO�Sa�U�a�b@�؏��FFI ��	��~���V��`}��w!f򈒒�Q ��Q��c��<���r"-������D�����gh�l�l�E���-*D��]oX*X;�T��>+Dܤi�����b�����VII}H/,�N�r����ZL1�b��T��%��ň��<>]&֯�HL[\HO�hG>�3"8���2엨;b��$������<m�;�:�AxZ���k;Y:Z;��;��B樬���K��ts>����Y�H|��}nbb�J�b|b)�#�%�i��k!bIП��I�>����|j(���}"ufz��m۩��JK(=p�u���E�ﶶ��/�êu����RRҟ�k���ϯn���~�8�OC)[\@��S�	::�(���x; Hi�}p��ڛ�X��=[�X����F���}�o�H����[0ر�����8�^���7�"&:�z�)��i��$2E}�%�;�K��WZ�����z��N Ŀ��#��w%6�Gf�!y\8�c���!/XS�d��x�������`v�M�O[:lSU�*!���H���q��x�檪�Y/\)()e����4�^�#��ߋ$P�D1���D��;%�������TO�KҪd��!�Ee*�L���.�==i[�o��?�=�<Q�-mę�-�T��2	2��l�ba��b�36�IY`���KGggyC���`_f���ST�����iNOO�{�߭���RM�||��L�N %��[f ��t&;���/.���,ªt���~٭�΄	J����~��V�K�c��n���� �V���m��"@�,Ihd���>��{�����A@���� ]W�'��t�+n��|Q�:�i ?������_}@���TQW�}_H�g��[ A�J� 0��v6Xgb�c0X��Oֺ0��g���!bV��u8�Z���ى>����X����*1�D4��´��3��Ŝ�S���?�j��>�D>C}�;��}�"�ڞ�c���t�K�ԭ d���qݞ��Lf�,/�r������BH���GEd�r�MO��b�Ixv�&ò�c?�q��u�E5�9+&'!���(��-G���e��%}�Z��(�������ӽ��)'		�\Ea�0b���~���[h륇f́��Ȉ��#]���b@aEluu�P�abN~��� 8����#������\=)z���+ͤ��^��'6��T�����·���g��HQ�q��Z���ك��K�)F���9�t�=G�4v�`{0�=TSscn�B3W�哩�|�,"ʤ:Z m1��T�VI%�����7�AJ�Q��t���G�N����խ`�`��W(�_��F���@GǷ ���P��\v[�ړ$�dԯ8q<��)��RaDu�f1��V___Dw��j%9uV��t�A�*kT�r�G���`��-����P����因Of�|���օxw98+��i�	��G7��i����m�=��B�3����ٮ�����4��%���Iin�t������h\�8⾏:����}�615�j2��P_};Ѳ��H����];�L��du��������a�I>�F$���<����@\m|9\���O�;�~6���snY]�اߎQ�P����#��<����^�J 9GG댟��j�$bq$��%��=V(j�6�"�Ey�=Z�C�>���'#��法�[��;���Qi�JR�RN�j��Q�չ���O�E��M�X��QM~���lmv�t�1�dgg��+���x(�>��=����p$nĵ9˺���S�֌�#�� rR�ߩQD��P��H�	b8 �E����U�<JQmd��̛�_"Fm@^��gr6B	���X=g\L�Îʷ��U�X���2oW갨7��߷0ӏ�	?��>
�"4����|q��?��{O�ϝ�ْ��$U<VT@�\JA���2&�#�C���.n�t��w�tX��oam7Ai��Dv���ˑK��;���'AAh�*�X7��ݤ GϪj�i�$v�{��˛	*<'gg��4�����p2��*j���**�!�!o��"�p��E�l.B�TTT"!��oλ��Z쨟������Ά~��{0��v,Ue\O�r�LD8�����Zg5^�	5�����z��1���鉸������@_��>������?	:�'^���Ǭe��Y6��z�N�Gm}x���dn���xX�r��@s�k~M�D:IvG���{g_�m�l�j�ơ}�"6���fb�Վ��f��p��K����g?�ݥ���2x����'�@&I�
9�*UQ*g�6�����-.��]�q��>���I�.�fu��h ���.���O�h����M��`�lm�]������z?/����S�Rut��y��͡b�u�E�q�n>se���2R�H�E�V~S������!Ǐ�a��,��9��lvo��Z�f\P	l��!ğV��&'R���L���.!����H�Ʀlm��9�ջ࠳y0��ҽ�8_���L�����&��!���o~�)�*! �x���, �BR������yV
����n�?a����މ3�Е6�AM�[\�=Ġƭ6��h9O��l�����x�!(;+����-�B�������7�z�@%�b�ؾ�H�ie�=ڡ��~�E����&�:�s��2)d!z��vK���2(�>z�(�ؐ�����1Pu�7ň��El����{���%\�J������U8.�>�{�����BG�]�i�䓔�U*"jO(_/�Y���#����������\�u��i��`�i��#�?l$�.K_R�����3��+��\��z�H�/A��*�D��a�Wј*%��˹y[ߞv4�NC�(-+�O��h�4]�7@�)_���4�xsc����1nΡW�2 �����_����5{������O��`4��v2%�����[Q�.B�bĞ��݃���g��o#�k�#�#�\� ���� G:8�>��z�I���e�A-�۷����s��.�n�p��)C��b�~I�\L��(�ņOCI�$���Uh"����,G؝���6���Ԁ����+�[i�~��&��T3�:0�¼�}Q���ijjjyW��7�WWW��>~��h�4�9���>4$+o��Ӄ�-�	�
nd��9p��\_͕,.���:��P�o��X?��:�o7��)TI���mn��]ù��MrEC�>�`K�������y�yj��n�6�&&&��s(��gp�\���XX����y|�՞��b�T��� }?�'��
�Gn�2ѓ��q7��sD���H6w�G�/]ﵬ�\V>i�|#�|��7�����/�G6���{��s�=}��>,6{������[��+>j��E���Rt��Q{ǿ���,,��aP�o����7rF'���R�Ǚ�P��?�����onm����x�g� /6d����@�F���W�1 1���.4�g���0�v� B;t���w�"rc��~��%�H����"}:7�������S�%&_̸FFG5��e��3�y�*D���@�מ�|���!s����������/�ٔ���
�d��4���C�Ie<�KBJ*[mh}у����m�~�����ȋ�z@E���p��d��J�u�����(�!v|�x�0HjDB�/�CT�"o����H��]�O�1J���,�b�]~�A�A�
u�E�H/]��Pw�?�������`1�f��my����	�ﴤ��U�d�����n-�)ii����:Zb���Ո�nz�<�&�&6.v%�Z���F��=Q-u-���ٙ�����S(G�Z��S!knׯ�V�p������8��04�$�z�`�B�w����bG����`��SJ,@	������c�f\��sa�[�eAO�#�7	c�R8kn�.`�#`;%l(����pI��ID�ܷN���b�����dq��T����{�'�B�m�Ǐ�?�IY�¢!>�KV�P �8�ʵ���t8���m>;��������/���W�)O��Օ�ii���K�n��m$�{hvw���Q`�j� �uK&�"]�y����`]j���0b"i�;j��li!/Y���(�b����]�f1�*++#����7F���֫���K,�P���vR>O7��hl��
�]u�$�K��1�!.&;;; �	�lo���X����9��z�	�֘̍���{�[��Ʊ$���'�9��^K'e	�`"}��*pD�)))=ls4�1�j{���� AM��x"�8Eu�0��;��]ي-����ܝ���(�̘9L������%�K'ʪ��J�X�����#.��%Lnf���/��j{�\��J������k�Z_�g�+�T�=�O�r��%��򐾽I�O\�ao�ϣ�	�*[V��e���oǺ��`z�������`�dHQ�63{��j�N2�w��Pm�zqDM���g�%%`g6|^�K�JH�#N���V�Kk ���Gszr�@�����e�X}�M��D-쾴)������Y$)��w��[[���!�p�`�y+@�VB4,k�|"�A��S33O�>�������Me���}�_62Ue��w@��
eHK#q1Sa���Z8"���ܺ��)w����;�����[����g}#�a�����2��Z�c=�ץ�Si\����خ�\U����e�o
Y�}��C"U⦪e�-!\��,��Q������5J1jj̜Y��1�ó���9��0�I����-�'¬�Td���Նw���^~�%G�u��M����9��E5�j^tԋ���,&娨��H��ݽ>�(d��jp�i�g�ͅh��Z��{'{�R'@�ԗ�ͫ�������@�����ee�_Q0�N��҆�N'1�yy}x��(n#^P	�O%���k�r��t���"�K�?��޳�U	q|@ݣ*{�$ŕ�{��t� 6��[S+!B"�/�.k��x��*�q����v�[�W�j�sݡ�����ar��H����������Br^nş�"++��t��2i�}���4�5==��𜊥��z�E��E�8)1q}����WQs,r��(;�
Y%�bWK������0'5��v��������%��Ź� ]ʖ��T/��]T�ME��j�<H���>d���֥��캖��K��B]�M^�K�����?���Ɠ��a��R�G�g����%2�O(+)Θ��l����z$ Kj���'��������e{@�ƴ0��N�g��agg���y0mtL�QR�m.B�'譳�
�k��G>85g��1͖A�T���O���������I��W,>U�N��3K ���.W~�|�LaR�%�HlP����cߔ_RBZ�y&v��GN�M���F�!5$/«�'�@�&t��yo}܆���> C��d�B=���qM[\־>v;��8��y%�	�¨�hn.QQW�74$3�h
Ɩ����m�G��"��sP��
c���ǂ� �&S`4s�5�	�m�mo�~[�L|g�,"2B.�}%���\5�����.�z���Ӱ����OV�.���ʲ>5��5r`M����fc�Qu���C06�T�c�ĒS���e���A�����g2�$�ϐ�t�o�'�1^ο�謾������K��9-v��V
��R�����ܫ������� �� �ozz�Z����􊮏���R���(�2:KFJZ����d�sƭ�D�)**�C��#7W��� |/�/��@�������<v^���br�}9S����Y�1�
�d9��?�bb�Z8挙����1C���NNp$ D�45D̪�i�s���% ��D�k�)<�}��2��^mX�&Ω�� �\L�O�k_|���}{N��+5�B���d�G�7�����c�Hn��wi�ga�ՙ<ҫ{6F#G'�p�ß�!�۱����2�(� ,�����?l�r��+��}��*u��D�����?B�`ܥ����R{Y��ō��G9/ V�|*�\OǚѰ�#D&w���3��#[��,rF����D�܉<~�?1����ۖ��P��V��U�i�$�-)�{���>��U}�azNN�ɐ��1���Qı������6�1�����5�_زDI��s�"=+�����?[^�Y��Y��H�K�_!�D���Hz��B�T�d����S�`Y�����=O�uJ��"�W&��߿�;���j��'P���J��n-��ݷ�删Iu�:A@���Ny��g���%��-�*���OS��>;�6�1RWoJ�i��qve4y{Cs*s�I���D�MC��X����DZq�b^�s������=���:%O���t�7��? u:X�a����+7�������QꏾQ�Z��@���޻�"��x����������n�=��ږT�+�c.�I
O<�r���MݎCI�^N �j,e�QH��)354+ ) Fh3ُ�V��E����a$�t̘�����}чoa^-�	*���1�/�5���V����H��Z׼�2H�
7����{�%����J�C��7RTЉT~���ih){j��ߍ���y­.��F���C�$O��c���s-P���Z���S%�̆�9� �X��.B�E�X ��?�bX���fY�W�iǒD���@�yr����g�{�߇���e�B@a9x�����$do\љ�DW�`.n]��rb�n��+���/{�eĩ���l��l��2���{>E����Cx�/����<�����_cPw�;J�����-| �Ǉ���6��,�@`�Ňz7���;��I"�0$(���Ud8�X6�Z�h^��RC=�u�<���+��@'�u4-m�4�"@��?Q*�I{S�����VSYX"r0-�I��ci����%��9�c�t,In�䗥J�{!g�������5\�h<�$F,�~�ܵ�(�8�m�L�N0�)w��_z�x�B$_5��y�;��V��K�r}����X�;�%.�_��ⲁ��kh+*�{)���>a�>6F�w�a�_&kΝ�y�g˳�-�dg�B'�k?�d��A[��o�C[��II��Þ}����@�.���~����?Yr98��S[�L��*�*��D��oH!ӛfa��rt�N�ʟH�(�#�B̶�.�R�}�r�jS*R
0����Mu#n"P{����uy����-**���Z���4�i0X����)��Zm訮^`X�;���!}�JE�᝞lo�'�p�
P
C�Š#�Uf3�
&�Eaǖ5��%]�F-홙2죛~p�he���g_�?X�������>��2���a��Vd:5}0�b������'��H�+;�q��9���%������G����%�=�����P�y�o�Qz��uL�**�}d�9 >�DEt߽���������[��ໝ?<��7��J�ZqK�.;{JJ�P'��X4�X����b;&�H�ŽoQq��˓A�ɇ�F2���L{x�l���V�|��K>>~���FΠi[t4a�ت��N�TE�N������-���Y����luZi˩q���i�z~a�-���fI���'^7��3����G_
t�a�����g9���Wr3�C�44��>�3&��I��$1FǑs��)�8ͥ��Hx�����ԫӚ�!'��������5(�x![s�X�[C� `a���9�<�{Q-'- �?(�W�:	;��L��ƣ��λ�S($ć����,J���A_���(�oR\܈X���N^�E���$�$ǲ�X�C�d����=%G��l��.�MQ@�g}�zd�K�6U�v���ه�MI��&�����3q9�������f�vR�AX��C,��WBB��K�)*Jf v���^ҫ׾Ŗ���������Ϊ�`gݒ.v��Ϙz./(����c7��p�(��[ �/v-�����B�3�Ža��o*ll$9p�+rٌi��-� ,�1X,O�.h�3��&��� DJJ*�2����u�����}�S@�#����z�����èZ��{���/��c���w�����q�A~X���_�튫P8 }rh{Vb�11e}��&�2�Tps�o(�2��6n�v�ݨ.>H����g��:jϏ���{7�ͮ���8q�6 ��_ù}�����s�ܜ
U�2K	mѴ�y�/�#�n��:v{�*q��_y���]X�CtJ��T���뜧���ɛ�s/���O}Y��W^~���m�l�59 ��ϣ��#�u�y-%�>#������t��:���_�xx}�l$J~�u�k	hÚ��u��zFNl��'2�C��.�(4:{4�~dt@b6��*֧=��s�I�Ð�C���շ��:yc_~�U+I5���8�����!�$I\TĔ
�2|P6YO��aX�(o[T�P\Yg��!�ǾO[rJv�ښ��C��Qι���b����8R�=� Y}�i�i}��C�49�����R�:T���0��M�iT�UY��A��߿�iLPBKW8-&m[�W��m״�sS*`��#�K�{�F��s�ǜ)+������E��o51����������&̒ȧL�|�%���u��P&�� ���N[y���t��T���Vm�q��##'8�k<��9ɷg�STTT��B����7�B��\à.����J�.7�r�rL1kncN�ڦ�ۺes�s8mG�\fqgE���ӥ��'T	rE�����>o��<�T��0�@g��}!H����-v�W6.4`�]`��ͅMU{����������BǏ�����~��>�"��m�Qf����]��.77W����z����&5��>�N�������a�^{��f%W+!��N��$$�E<4���f5�z�'
8��P�7o �e7Կ�Cp�s��40�82
B��C��&d�����f��A����)]Z���-Z���D?��:�lW�����+������_]�<�4J��IR�X4��iBJX^���s`ȂqG�����"����C�[�E�}�� �����!�����%�C����������H9"H
-��0t>���|���p�Ή}�^k�}ֆb��D�����UW��tq��y�gkmy���-�t�Z��� ��+�R"��Q�wm��ٵ�=���5�nT`��gzU���rCC�l�D������`s{S$}6��jdf��'�}�L�5Bش@�᝵*rfq�nH2>d�Y^f��֭��OF4����Yͣ�
���:�!�8�o��g�����w15=�z8IH��'x	���jji����uo<kI͆D�lhd� ��'DWN�����{�A����՟0u����'+��M��y��� ��tv�]A�]{��*zi�B��ǆ�����,�����=#����b��T�Ǩ��RƷ<(e�0aK==qZ2Ҹb�܏���S݂Ъ�f��پ�Ñכή�ڊb��!s��XG����ӧ#[�w7�?�blu18H,$�p}��5d��\\\�Ƿ�N%��L7�H�l���v����dwf��S>��XJ�l���x��C��GHXȠsƆy]��|����s���%�I�6���'���R�ă���E�� �`s�M`c��� c,l�$f7�y��^PB�3�P�V�)����Q
��I]���a��eb`�N������g�z�{s]��3y��W9����{�Z�~�K�E�4�PY&���8G>%ǫN���G�&�f&0(��[l �Ʈ=Ykɦ�,�ذC��Qi��w'��H�i�����M�D��(�V�a����fP�"[�h}��_�T�%�{�XX���R��eܙ�1A�o����ׂ���{=��W���l���W���3�D�o�j����?���0*��4U���T�Ǐ�-�TcJ�/4�}��&���5�/<�̊VZ��=�䉈������ei�$YD�cvan�p��t�֛�J��I�����w���i��G�G�dsҭ�Z�v�/�j�J$c��I�XCD��;�
Pa��� �	���$�bd�wN�D�-���V�`�bqj��'-��7Y~V�h��Z�r��6:q��r[͇C��fd�����W~����mI��`Ld첳��#��!�g�а�C���*k��a�lz\�"+&�&`�O�'`z&틭\U��J�p�����8ȳ��'f�lȋy���pX�=�A�U[w��9l�qN���ݳ]�_O5D�^h���)g����i�c�B�t�] 6��m�9�h3C���e�;�������L�?�0)	�84��{Kpbr�؜��8�(d-���~�9X�]�Jpp��h���4Z�C��fhox�W�F漲�?9N�}g?k�5G2�,�r�ւM%�\�s��fng�����UX�̻ʛ���q�'�����WT�������7�b_|��u���I}�Z�F�u������=�tF�֞x���?�.8�l���",�7���v9�[C=E��~Y�
���OXXN�}}J�-���($�(m�!൹s�$"�}�)� $
hC�vQ"��ԣvs~G)���Ɔ�+��u��~���q������Ĝ\\�z�J&�*��D"��ފ��F�0꠽E<�*{aj�~T�G��`?�	�,L���ȐyA�UA��1<b���������=���q��Z��R��(�����_�M�y6��ȥ���Ӽ�q��|z��a���kI~��ۉ��YVf�$��1YY�۳�V���p7�W����/e�	Rd.�W�h�� �]�g����k�����iv���W�|k�UV*S�e/_�?�y�Zz{̄��!���~^N�c�4�����h�~;�N�|�Ug�B��dػ�ߙk�Y����!aӟ?��/�YS^��b���%�"�%�+x�p�G�]��R���^���f%�%��t�]��,��g���e�T!K���=(4��W2/���V6b�_ZJ �b��v�1�.	�!�Wll����B�H&��A�]��$��j~���#
TX8�i�y�*�,�Jz��J���c�@���^a������M�{�u�%'���.9���~}}�n47 �O�Je}B�����T.usJ=���������f�G�q7���Sx}���iσ�Q�����m����ED�?['Ο3�Ⱦux!����y�<�~��Z�������>B��yk/NQ?���˓�{�ٳg�����R��A�r��鰿wl ��AR2���T^ޮ����9K�h:��EOl��Tk��۱"C6ܹ��rZ[�h+�{�Q�.i��phտ��؃��q~Թ��<�N�'� ��&3Grѐ[� &i����MN�j,���/�Je:�vŁN"k\8���0�zhju�]���*����mM�s6))��&����"C'�Mo�U(B�@s��k�3�[tv����sP��Qd��H�~�*�8 ���o�dy\��Kp���1$������zP���&'+��������ͤ�@�﨨6_a�o�(��wI.�F͘E��h���H^�?7��^<������� _�a���f�]З���> 0�i),z#tJ��6�/7W����'ff�M?ME�1p�{ �KDD�I^�QO����J���T}v����������`z�+9��?��;T��}����Z��fq:>���U�"����i �<�y ��I�l�NO�]
/4�!���L�߬3'6���;�-sE@b?�el���MR�O�D�旙A�����"b��I�{��&�8EfsoS�?3�eX���A�­\�6�ǃ�~�����Zt���~@1`�V��y�`�}qE��KK�C6�C���v���<	]oz*��É�t͡� �EaҢ�W��Q�ۼ�8P��F�[�Ĥ��V���ťBc��"��1����F�O��
jk��9,Yc���צ��7����e]( �C=w\ �G2�&z�`�	�]̙_M)�_
�bl���=�r�����A���b=)��yvߚxy��&�h���ޞ�[��{	���/�	$9 d��CC���;<W�vG�^�����qZPP���."|R#�z{zeE�P���x�q�}2�Fсm�������/�{y��DXIԮ�=�=*��P�h!&>��\��% @.�����3x~��_�m�H&�A2����),d$.���Q�z�)� ��r�оD�8y�(��fܭ5Èc����]I��N#H2W��n���q�����G����iy9�r�M�~d��E�*��1&(R��Dcyŏ�j�CT�七`��Y����֕M�|e��#�����Ts��g�G ���tvNV�G_$����е]��G9��Z@�l�6�uT���FSg�f O��`c��������!yd��n�g��IG��	jF�x�oLw�+jy{
��1.u7�������Q�1��$��k�,��~0��m��]\�ρW4���2�
�:?66�0��-%� �FwHj�R*�����;��T`o�1nd�����!���~X����������m	��; ���	�~H?�I��������Y�:*8E��!�%]^�5��|��-�~���~��sS3�!��Rh�%S�H�����cu�9[�\�D���	�� �>�����v�]���>�m`]q�QAńX�-�����4��Qqa�����呅��[���/-�j��4zzz���/��s}
�c$��a���>:0yby9���Y=s~���v4�
����B��l|�Ρi�c���YTYIQ�$�>T�b��zХ69c��,jF=%�2׼�jv!b�;�!"H�GY� �W�.� �$$'���A���^����`��X��:�Ѹ9�<+D)�E�Ş"eUd��'�$�ʆ��+~�P|բ�f�����8��۹8x��)(�C|Pp�D�Rx�Us�gOu�|�	���G�h,�9�Eon�S'qr.�dߊ�'�,Z�M��������p��d�t��/��4O������	���/���6�`�p�"��	�^Wr5�RV|N�K7�<�w��dJo�\�������f\�H˛#  �}3G92��5�ņ�zk+rs�d��T���;�بP3U��C�ΚF�bɯa<�#�$��	���⑉G�=�i"4����u� o1Ek|�[7\2�5j�¦o�}���ѷ�⌄H�}��-�~O}*c˾�fm�� ::>��D�����SM���I7>n��?�]���a����}��L��s��j%��݉Ty擨"#�ش���ٴ�`,>`�vd	��L������*�P:��r�t䎴�\�d�Cy�Q������>$棇O97��������L%�����l��;d�>��/��=3-��k�B�x�r�LC�Q!��K,q9�k"���P����b��S���ٌ����k=&�������v�&E'�y����V���$oѭ�
���}���9?�R�56~1�-�qj4}�ϋ�*4�Ҟ�w%}�������c�g�ޓ�� r5yi�;h,H Mڮ�哯.><���.��.[�r�� >��w�6
�5��&��I�����.���Ռ+}��'�6*���c[i�lzQb�\^O�Z�q��������2a��J%T�`�ӏ��1�m��u�v���pz�e�.�9�K�+��e�F���BΑ���#~n�i���a��I���^�1�����~���Q�I�f�`����p�S ���?:*631-(���%�\VV֕L/��Q<��Yc7�=�P����?T�(�ϰ��"��-�䶔��ӳHI�J@ˀ�~������z�
j�`545��=�M��9%�*ʾ9OAmh�T�c~��n��q�~~4X7oq���j<����c�j��-qx�����x%�!�:���3���O��IIK3g<��N�����O������PY2Cث�Jb{��L������N+R�g�K�0u��Zb�7���S}���M����h��ZH��B���ϋ�$�ML�	-4�U�f'���
>}��b��JmN�AS�t͸�5���e�5���������HJ��Q���/o���0�Q�O���=��Ԭ��� ���K�Hu{&�MV�r�45##��S�<��r�n��Z�[�/{�⪫	��������n���õp�3<�Ҫũ3�p��x��G�O���p��a��<�N�꘽���n�>g7�n��i�PCOj?�p3
X_C-��%ǉ�'�[��F�ۍ�?*��c�xa[�����T�w?G��/�?���`Qe�yn���M>����`�#P3�G��G����= �W�EiZ�ā����S��V%�8lJW�r�C\�98Jp���S��$9Lw'�G<x�!i݊,��삠�L�$R�찞á*zP�����%����TpI�o��݃�4Z ���N�$�`���i)A�G�z=ݼ�}�E%��q���Z��UX��se$d�+GJ�����Js�����a�j���3L{��:8�i��U�[��o'`�2�έ?	}+�� ��d��~���N<ؿ�f��鍧Z>�cs�_NCx��S]��*����Kek�Lg�W@ �R�	�B��T"��yz��a]�����m�0D8/m��}���ߜ^�����Ϗ��0H�����éȉs*�U�=���̧��r^���٥��芁�HH*9 �8��=�bZTP>��F�'�5�N3���(5�^X����fdS�0�-l�	'�-�r͝���^��w���?[�cH���%�^��7ո�{����_����?�sw�V�}{�|����oZ���	�����S0�{��_�g�`�K�%�	bu==׹��T�3��s3H---C�c��V��@����3)�wv��z��)ԐE_��蛘�5��|�/��u�7�,siVB�dL�`�{�j	��Ɲ�d�~�&�{GJ&&O}^�	v��SA�(uz���qn믗���uG�_-Kb&�V��D^�뻖Q5�1�UW��]A[o�_���]�,��3�Zy̪��#�Ѻ����-���)���F�'�b��1���`�}�i�����ЊR���C�S��O��jj@�b͒@��L����+�QR�Wnq2O�:8�;�������m��p�H�:Ϟ)mVc�M*5Ya��=����t%^{���x��m����<Ӝ`G)���~-6#������4�K�n�.���d�uLR�Qn�箲F퉵ނ�g��䧟85�����mU�&��T�=v��Z�r�rޗ�bm�;���M�5����-r7�๿BBB#�Qs;=���&!�W�{+�+�s}�ʌ��3_�چ��C��:t�(~��UL���ߦ���-q:��ך�g��l�1Ş�4�W���sX�����{�c+� ��$俷(+s��~K*��T^�{c+p��@���@�p�9o�1�<�.$q��{#��!'$_B� � ����DNh ��Ѕ+'��g�u�戝��׮g�"���}0�X�C�����U ���Ş`R���l��!!!��h+;	��<?�H��]�c1�������mw!T�
�7�Q�}��I���b��ڧ�w��}J�6�@�! �:iK��{�6��c>w#��Uͣ�H�m���c���쐿��O��X+�x��ۅ��AKm��{�p��r��@=�ŭ�Ü��=�i5U`��2�^����]	d�+�""��б#)�c}tsD��oM�B���Y8�D{���H����td,xV&alm5�TٌK�G9)�ɚ�ӷ�3����m�K���ȶ����g���)́��Z��G�?�yN/1Ù��z��:ů�68��i	$T� �8���3����	�>�ȁ��[���q�4=fiƀ�|iM�����?��9��{z��8^��5����_+*�!NM<]JJ�`w�~	^_l	�ZV�Y�<2 ��g��r��\`"���򟊲Jg涭Q�rt؄O�1�]��]�{��n�����n���|�η+��a7_����f�QM-D���9��/s�C)Kۥ��F���_S7��cs]�³��?��YH�P�~|��7��Xb�����&���L�ߪ�"x����P�el���-i���6��	Ѯ�pN���-�C77�_���p�B����P\
�e!Y��:�{ȃ�A�/�Qe�������nQ�]�V:��
b������w��{t�t�k ��//w�R30�L�JL�l��prm��w�Pwr`��m�wvJ�c��׃/�z-������n����!a�H&�]��IY���a�V5j��U�lSnB����f���a��#� �
��7�K9��߿9�ڿڌA�$d^������V�a�/����D�^��1���=h�i��0r���Gj�AQ�V5�t��Hz��s0��]d��I��t�I2	ö��i~Cn6ٍ���Yͨ{p��bJuu����n�[������I͓���%*>9�(�X��;�T��Z�N!R�<;{��)���VXx�i ��.�f�d��vsw��.�zv$q���Te�fka*e�O�m��U��;ն`��sM�x��0�SL����������Z�ppp�..���g��
�>��,�"����uH�[�Vh��xqіN�.<��הg���g@�z����ƙ�h_q#3T�T8��5�u��,l{ ���H}���w_����f�Gu�Q�.Y���A4`y������8##}eT�1δ�)
�$�_f���N�0��=7f8�b��t<�ZA�2�Mb~�!k�W�옩�d6�wC�%��ׯ�d�p3?����������/����#״͖Dd$8���bQ���|b���ӧ�8�&[ZT��w��␱�Fgw�H��� �����~�mv�@S�?~��LCysp��O�g�g-䥱n�;NŞ���h�L2ɭP~���',hsc�vX���;Y�(g2��T�]i��< c�N��0�}Ep14�B�� �G��?Q3�w����B��c}{;��/
A��+�I�r
L�A``���g��P+i�U��dy�WJP�@� ��R�oP�AS	ج�8��T�9�cM���HV���V�@ot���V�mG�|�J|���K9�:z�Gu��jk	�����ȷh�jvu�q�u�H�6���*����кt����$A�l#҅[c��bK�8.�fZ�����B��ܕb��c���i}�ߩz��CL�sp<^,��h럷V���A^@���,���qN�5,yw���{ʂ5:�ptKaq� ��}$%s���p+|c�L"�������ru���1�U
^�	��fju*ψ�X�Wxd+x�x��UQ�Y^j<Kff&'WOQJ��N'��aQ�����Dʜ��VK��Dl�qB�Ftz��I�����<k��Y��N�~����� ��/%��S�G#F���c�I����Q�Q��]��	��P'�~���Z���fe�5oNW�~�E����i������\���2Pe�����K����_��8�C7�F��>ù�ݹӧ��7��&��na��籠��v�Ĳﺢ��)���-dj�z��{��ӾtM�<e쟱��c���N��6tb��i/�}�,�[Y�"OVZ��4���zK�����1̄�r��A��� ���R<x�fΧ��Ń�����0��{W	x������.�=\��\��2r��v7�T�z(�gm�������zs���af��ECCCmD�������¨WD��팖�r��	�PH�/%y�V��ۚ�g|K��H0ã�����GC���dq��"�P��
_��JO�ˆΫ�P��ў�}�n���'�uh�W<�3/�ü���p��P���������
Q ���TL��% ��yy���V>A7��T({�C��o8f�qX��Iq|̓�y�k�n���cn(�e�HZ�wv���̭͗��15����� �I�����2kE�~�Z��7�pA�ZӰ3��ҬZmd�X�����,D7����Jı���JQdxWu�ڇ�o��C^/��(<o<���e^oЎ�mi�g�#�+0�P!���%iz���wXX���;�wV�8�QŚI2�n��ݿ~=���dkn$�L�f����8:8`s7�h�HY�H�)^0�"麻�n�+��Z7G��3^m���X1�̞{,����]��C:�Wwzq�������|}nAi�D�G�|ɬ	ݎ����s�ߑg ظ��=���I�W��\x���hxX����F3�M���@����y7Xb�<m_9�E�0��{��4JU2/�]}�qI�#��-�[#=������g��O(�R�k��؃�� I�E�ց�<�rp�L[O'p�R���������͖<��[Km�����{z�w�5��r��IW�i�-_��c	HWr��o��� ��a��΀yf�4��"x���󭷹߷���FF߃�`�=j;E�m�{:`�tt�ґ�?z������������,���xǏO���a��׉��'-!����^���A��߷�����!�[����n*V��<�d����*+ô;f���2:�ȡ7cBr�#��8	:�����9�l��v]�L����a��/ϷTH)����#��>~���4��[�91���d�R|iy*��ЎHP%�2	#�nl�d�g ��㋫VdBڠ���EQ��߽|�dk!��ef��l>A�� Ŋ~���U�`�,-i~J6.�J7Omu?�4�^��՝063�[���)���U�4��XS��������{���Ù�p�ݐa0��ݯ~�|���9�.���w��?}��*_T�3�aڷ�{ۚYes;q�vq��Y�:.P|Dӱ���{w"�M�&++������ɻ��r35v5�r�}ILk,�!TX��)�KK���:��oMU��8����N��mEƫ�����ۋ����_��H��Y3��<����y��Ba ����#\�y��%����ڹ�o�eG��o�:��{�Ⱔ��?a���#����:�$0M�e�5Jv�2I��4]���Rkt*�"���4��l��U;�k�|��e�G�
��O�9�����M��������@�K���%q����+�Ļ�焄�����+բԌ��������D������(o+������`�d�%H�g�C4��\��Z&����`����D�U��@�,�p"$d��;�-t�����^>�N��E�m�'<D�O"o̠>� ��9'�:.w�v��O�x#۱���dz�8�Um���'� K�n4kn㎱P	�K!���nri��Nh[����eqI�J�P6µ��p�����b�yg�ƚk%���m^rB��0���O�
�`�����;��="ïC*w�U«x^��e�f��ukv���{����A� �32�r��*%Ĺ~�P�Mz4��E�%��-S��(Q��Wyj0���F�KLލvp3�0]��k���9�˔fD����d3P�D�!&��ب�)�����~J���@J����}�����O�^���H��SN���2� �?�#&!��X����l��l8R񾼏br���%.�Q����L�6tGt1�gUҬ��:&.7Ǒ}�'ig��`����&~�.��vS�f&+�SMJӎ� �DY!#c�w0���������۵��G��Z֑�p�vq��#��z�l�ͣj4���I* e'
F���S�h:r����ׄ<�]���dZ������q)%z�������tϞAR�aD�x���Ox�����JJJ�||*��8!"x��`�㈒�0r`S�K�T�]T�j�⽣�7>��Ѽ�u���.��h�܆�R՘�UF�$����U�К�KK>A���<Zi�ƈ��o޼���1�.I5��:�)�S�R?�o`С��J���=]��C~B �+$,���K�Q�b��ء�h�ѩ(X��C� �L��LЬ�C�=��U�	�(6���	�^���T��#�K��>��`��fF^Q�|�hLǄ}!�tn�͎o$U���?��iu�G�L�j`��;M�	n�Iq�C�8ſ�6 �>;	�S�ԏ�k! E?66n`b���]1�#;�����ZԼ�i�F���j��1�պ�*	[� X�5��PS �:�4�))tk��_��M��ψ�fҗ_p���d6�Kz�e�-����i��Xz>�/�^<��+���"�utD9�����7����$�sD� ��������̷?666)�/����Hp��21���oT7�h���B�֟�?C��h W߮�͊IR.3�jnm��%r$%�@sW����G��]v���2�''V/1��������A�U�<x�V��Ve���Rf^XL]�v�iT�A�����o������@����4�����/&��'���|�˨w��.�Q�H[\4�U_�z�*,ة´���"�����#Y4�׶T�զ���+����D�<�,c#.j?x� ��@ë�������Ui�L,�����pd�e�����	@\��"vΟ������ߞi���\،K���ՠ���X�:/��a�Uh�4;;;��~rB2o�� �|��>J��%�Ww���7� ���*�ֿ��$[g�sA�nT��X:�v�ׄ�����.Ů�L��4�&vǘ�3�3{ST�W��̉�����{P�9����|�������D�g��F�������6s[�_��q&*{��qq6rOE=���f�5֪#�����x4:[�gJ�~k񴅁A�`���h�=����k=]2$��qGٚ���_w���"CV;�r{��~0�l���#n��)5}�
/�1�����9v�P
`i�v`9�L������d��V��V!���&K��/��L�9�5��'U�0K�)_ΡήO��c��*�;{푸S�6�M-�����&=�2/���ޟ.	A--4��������INAU7���ln� �5]����rfg�Џ�0�︞|a�����647;-�u�].U�p�r�ȳQ�DW�pO��X����
������U~*=@����%�1�5Z�i����F��?���ha��g����	��k�5�r��r���l?~ˑ[	��z�|R�E�}m�QĂ ���ւ�C���<�W=;�35�kP������"Ԧ*z��h��y��x��S�3���h��@�5��Uvfܡ���ȥ���}|�DB�_x��Bb��u?�]y�WĘ�H���� �1��ؚS������oH��okm�t��C���N��Y!���ufg�:ޙ�8��?�N���5h=��J��D+���=���a�_t���Q���`����\��Mx�����x6
/ ?��EĻ�I[��'����H�p���|����7em`ܮs'0��krrR���ڲ��9(acws����� @����J��
^���0� y'(L<[��S3��[�@�I� ��SY<b�c�"n��i3bf狫��C4��m��z�x�uH�{f֚�ʂ���-{�Y��|k�0"��� ������<5T�����������xt��xQ��US�0�e���fJKK�n
m�-��%*œ�����C���;Z���8�*n}�F|_����/_n
�Lp}���K�5�Ij=V�h~�w�dQ ^�!D��.*��7;y�H�7b%}����|�3�+�xQY|f���O��U�/�g1V}�?�%0.��8Y�m�tԓre[pq�2���3]��:��'[���=��[{�Gx��%����$�u���{_�%W�p���ʱˎ���sjr�}��cK�ʕN��V�Ѓ���1��$���j�I������z��zt����࿚�5���^�pw��z�W"�a�l��N��3�G��)?y��2)�!v;cd�nM����L_C���&��YYeY��Ϧ$�*a�$��w��w�R������%8��Xd���˔IE�����t��h�p]�Ң���o��ϴ: �|}�XI	��<;�BXUUU2e�6�c�����U�w��雡R�/�2�m��h�ڧRv|�J;%�^qM[Z�-�\��(��+�Q7�M���� @�+x�JxQK?��k�kNbI�8�=
Z�P�x\,uXIAU��qS�	B������~1����}1�`�P�Vn��o;�m��A>>��>��y��$^�� �9�Q�}��j�5]}�� �����t���p*4$�!�3t�;�ʟ?)���e�������ȷ�n�r7j���P/8r�//e�ڿ���"C���5���U�P���1R��j2(����:^��F���٘����T��`?
����#����@�l�aoh���7@�NfM��s>��|�+�VJ��v��E����Z(�o�z�.	�7�/��GCw���$�p��~-������t;�q�}S� ��PQ�tYI��
��k���^��� ^vz�8*�,@@�;2��ʠϑKAo=����;dS6��}V�4�o¹�X/�����-�"�`�CvB
8d��f�Id��.�~y�\�Vd088�7�>?��qY��[뉈�x��F��� u��2SV��Ӄ�����水���qp��O��mY�U6�ǏU;TM�4ȹLa98��'жW����o��`���5�>���?!(�;�}�
��h�	����ʳY�a^���-�Wv[��扳�í)��6�r��o�ǘ�=��`M���G�gH8��|LS 0�������W���X6%b+���c �4���c�e���91 ^�RJw9�~d��\L���S�	�M�� ��;4�2�4�R��p�E�E��t��滺pI��b1]G.�^�q�r��.��Eo�M�H,""r���T\*|J$������˧�VL���ɢ�}�9d�I�T��˝�	���>�}��w(jɑ����ՇTY��6�C�GG�3�<}��lV���ӶH�g��ͷ%YS�X�������徊}E��cX�}�ާ����M-��_�0��u�s���8I���1$v���H~��#<b*}pp�;/ɋ{9�n��ߥ�>�2I���X�e]1�,���(��n}�����i�M��_�HWk�<���3g��2h�����g��$6^*@�줛�Di-���>�h��������-������=Z�-�UY�;�a$�h����ޙ��V�n��M�P������֟��K����111�M�����OY���9@���//�vvu�V���0�{V�DY�Gӈ������A'zu5��ӧ%}S��d�(_ E������jUSSJB³E��V����#��*����ƫh`I^�$��⾺ 7!CL�.�2�A�J��cN��o��t�B�J?�Z&���-u���NJE�T���+��|����w�!��1���R#��S�^�l����D��wL�������}GC�C.J�uD?	�BR���'��>�hp�K���3�CO垬v6S���+��a��|�N����q�sc�0,����?~��8~���[�nm�[�װ����8�����P
g�����=���Ϗ�yW�!y'Tp{szDٹ�a�Bw�1]���~��1�ȋX��������L�����D�M=j�
uuv.,�^!:�f^K��+�l�?]ׯ���s/��s���U�/��j��]\\K^AO��������./�����!��؃�b�ڲdpom�5��c޳]���$F��+Q�j4Ns���l���[���S]���(v�хŐ���WP�Jy3��Rďh��ʼ�$���*�6����<s��)A��[7e\�mM�����*��ҏA���;�����[,��OQ��a�r�(׏�#���� � �r��&Eq���[X$4/EX>��
E	�bBR6�݃��v��ř���,A-~-6��Zv�y���"1��a��8�X��dC6I)��2���@�Ժp�;�G���#*K��Y��8�^�,t���1b�x� ���Cv�.�3�G�Ѡbz)%�xfnn��9%Uq$l�ۧ�
O�����a_ߪ�
��7�$w
s�,n�,��Rr�$ !~-����B��%l����dOK�{N�ڈ�+��D�Ycx�;��U.����ʠ���M�U�UA<�"�]>j}��!�%G��NS�����g���O���Ӟ���lȂ�fgf��w����K��L;�99���G��I���Y�2����I4�f8W�+��%M$KAu�����+M�6�h,��\	T�������-��{���y��#԰���}�f`��8Q�)�鄄%��ǍR ˝^�&���UH39!+5I�r��Ȝ��]2���N�N/���RX�D���;B�a��U��#$�<�z!�Gx����w�̿�ӕ�|��(��@;���w;K.1��tBc���)�؂�U6f�N�b��xU�`ҥ̘��Ըvg�3����_)���T�?4Uvv�S%V�S\I��ݩ��:��L�N�ZW飢c��o���M��ٿ�wm���k�YPv��o�-Usp�����Iz��G^q_B��u~ݐPL��;�(^):r**Vaa#�Ս��L��8?�� VK�J���[�ʖn��D��Y݃7��#!��q�sO
��)U��z�_��]���-,=��B� 
S�(y8��*+kc؁�57�U��[��Cnv�t߼�ע�,D�\�v%�y�iӂ�Hs����.����z����O`�k���<�.NxN�
���K`{4���R��\�b�F_ɶ�Ժ6#��1Щ�.�ee��?տ-E)9�!�q~�5T���+�������V^@`� ܾ�����M18$󂬩�sꔲ�nf[`�'d#)%-ņf���!( ��-�ɁYʆF�U'v���o[G�&.�H��Ģ"־(�m��A�9/�X��S:��⏏5�hS�<�!������CS��.�k�z�5Y�-��c>�s�{������N�Bh���#=N�#��bj��ܸ\T����N+�4S5�"=11��Κ	r�W�{��%i��jr���=�Z2�kiAQ���xb����o!r�O���r.)��7:s�w�[V�7$�y�R{���w����9+�YY1���EO���^��+/+!@Q�_���,<\zP33�ƪ������B}�dA�Q>OOؤ0�ʪ� �Bco:xA��e�X����_`��Ψ��F��P���&\�G�y���-�Nr�Z�w���Z��4I���qx)��I�딈	
FA�ne�0]����[����7�ւ� L߻����¢8dE�8�UV� �����"x�<����I ��d���*�_��u`��~1�V��xhҁ�^1xhU5���-���б��0��G98�P0��a�
��h{e� +����٪iW�(Y���Q����LR��̭�)_��"�]Xp�vS���mKII#vv��9�Pޞ7g�y��I�����׀M��r��Xھ<l�GaY���o䘝�-��)F7n���Ÿ,��ŧbd+��8e����	�"�jcx��iX�0����I���rl����F
޲� ���s��'�AQ���'Z��_a1��dj%�?��B[ZL����.�M����PRQ�g�c���/1����w� �2���&9�Gna�3#�:��GUUߣǗ��Pe��\�x����X�����/��
\Z�H �>E�׾
a�����l�445
q��[S?�Q�8ȱ�p'��fb�?Q�ȯW���R�j�eeu�y�sr|��ʝs��pDS�k�f{9��A|��,sz���;[�])��Ӗ�[S*��X�cqp��ψ��#
�M���$o.�G��xLk�_7L��;��7�`��q�SlO���<g�k8�T�����
a�m�]��-��l����rW�w��<���Ce.��wk"��@�����W��e�Ψ������br�����o���f�+���ć`Ն�u�H��o��p���T���0���â�5JC [mmi�������8*&���H;;	�����6ƣ��g^��O��%�!���=�yj�O'-����T���c��v��a��(�n����1����ݹ��?E��첉��|��!�zfq3\�T�m7�ZJ�OO�Q?X�=��+��H�	l�����(��m�\�CI�%�n�n�c�X�DDrED��[�[@@��eY���g}���]��O�9sf�{Μ��>���aSC���ɒn�\H�/��wu(��*k&��N~��c����;wD�����"��(�3��#'0o��q��7X��vd=6 ��yO��t\�c1��>0����X��nR��!�^��Gf���d���Z�mm�U돟./e��P���z��~�}�#.�7{��K��>�-�g��ɴ�hG0��s��Kq��}|�mNJ?�ˑF��#�E�����e$>(avF!#'~�,�|��k��z����n����²)�{{�rݹ<�;��⻺��y��Kp1ů��J?,��㽷z<�W�e��>�ّ��N�Z�Q(�����1������߿ԐPO�`1=���,[x���-^-�-�������H5;�|R�*Z͹	L$E����߅`��ֹ����9ީ9�m����]UQ�)�>������l}��u��&*�qd�kɛ��Ȅ�D�f6�6��R%�UC�V�锄]����u)�Wʫ����?iM��S]O/�������E�.�&o�iyTb�j��dy�(hU���W��]�%�X
^�T�k�����|-/dZQ��\��7�Wu�������}�T:@�߬��q����|�N��m/O<��� ��Z��D<�� ���F��(��pS;c�g�Y^\)��gQ!�>�J>�I���h��<=X�\f��I���o���i�����IDx�k %��1ү�c�6[ax���,I���A�C�Qm�B�VIhQ�� ��-���<I"�_[}�6k�_E������` �V�4�$��]��YN?*���R�K��
�dn��[1Q=�&�ȱ��`P|�h�Ĉ"������=|2~⋿�p�WX뫈�*�k�ь|��Z��;��g��g��A�7��E=���Âe�XP����U�3�E@�	��~�#G��|2��(�(�jX�� �}y#r왵�R8���B}>	j>��#��']_��Ҋ�����`����rV{�ɊGg���;���sB��$�xu�u ��F����Σ������6���<ǡ�Tbbbx�nq��vzŪ����^�qs��ng��C�g�.���|�kP�\���+ϧIV�W3MgZڱ�1H��-����@DW�3U�k�8	���Y�~F-���8|�'?���܋\[@�^K@[h�_�T�l�كB�hec33���W�!i���G\$v��U?+&��c,�Z�����)A6�''_�<d�_h@��ۉ�����h��%cJd҃�?=������Iy��E����8��\�'E-�����$��p��G�����+2$!���V6��3-��`J�px9,�%���٩�)��F��.�޸���lYj�lO�0\I��h����$o��8%��F�T����S�1k��?"�t�P8����mJ�)�"'"��0n���kX����z��d�ejmM����{�Su��0���_y�� �6���@���IYф�y%�>�EKD�~\.=9�T�=|H6�� ���������,��	���y<�9��yH���� (��P �'�4k�t��q��� ��TJ&*.�[���2g���/Ƚ��|&_��,�[b���`�#�o��gy�o�fq5�v�K��L�M|d.�xυ)Mh;��*N�dJ��<4���äzĪ��	�	b�2�;ۉ2��7��\��ω���\�	[�qY����3�8�3�H��S��ӂ����gHBz�E��͂[d[��Q(T��{��S�:��~��
�7D���s�h�8ylʣ{2���M|НE��?Դ�o����Q�SA�u��/��w����()� N��^������s�ѧO����sҷ���eY�ұ���{E^A3��a�k�
"]b���(V��5/O�BbUN���Z�zz� �NtuR���ph�m�x�K�,�J),�{Q���O62�/0c����EN�s��-cny��*�,h�g�y�Q�5E뫀�����9BT�sH;|g?0װ��� �hpI�I����[�Ō���;�1��_��ɷ�6���-� ��P����a�_����V_s��M�Ol��W����} ���v��!&�V�=�]�����j�sN1����c��ҡȽ[��ˌ����,v��[��<4��1��i)�|V���VBX,���B^�%��($֢G|�{�0���=����N�K����B׾=�G����$�z�JFųt��Hn:��v0_�{"#����5�y������Mϐ�)��m"���y�NЭ�ߪL�`�km@�|��f�_-��
].H��ٺ~�z��J1��r�����`��uP6g�$ɵ�xY�";U��G\���8z�6��1���"�?Y�\A������Hg,�j�����k�o�17>h]~��e��� ��~j_}��S��0���?x&$��M�����?�h_3_@[��Q�n����i+��N�/��#�p�����cl�4ң��z&��fF�ݦ,�������6�mkK?��v��U1�5׃[296f`���?��}|"��F�Bv�O�ep`����H�������K���Ƃ���}�gb��EM׿��.fqOGwq����z�R�?�	9����]����q��֙J��[����#	ڑY`�R`���$�^�#''�̀�n���ruZ�{'z����3Z:��.�b�̺���$H�ln��:��r>�A�d��N�T!�d�! ��hp+��Y�f��}��{���
6��g���Y��r�V5L��-�����5S��aMQs7� +�W���x?t�W��k��:iӿ񲬈��G8D7�g2s����Վ���TAs���9@g@��Ύ��UZPc�-};����"�7q+�
,�����i��Ī��s���L�s<�Hc��e �T��p�r���a��8�qD���Q*�ug�n�aR)�~����d�����	��lw�Y��
��_*c ��
�O�Ǟ����[d�F����v���`��c&��te9��5#v�֮���TG\����[����ȉ�#k��ggs_������{6��y�;�\���(��q��'��8M<���C�P�l�V��3~����D���P�Ӯ�<dY�YK+7vt�S����NN>"�B�)���p�!'�f��tA�E����FTA���������Z�33��]_Q�~�W��nՅ��0Vւ���e�$t��S�п���8&����Mqf��vh���W������Wjncc�^inPM]C��Th��q!���0��� ���9Tq���HCw�mf����z��}t�m��H$���"�_�p�������@(�r*Ϟ�Ĩf�5�$V�w&3o32�����M�����
Ð�a.Ԏ�e<�{��b.]�.[�*..���AL7��\�Ť�ng��b�.�)�͝�>�^���E��d?���$��qb�#�k�%�A���Ƙ�~7�H�� ×�ӗ�a������Z�T�)3&���I����J�M��Wx��r��Z��	 �AG_�������gk���=��	��c��Ý?~�
&0���D���?���k��4��v��였���+��������`����"z�g:�-��%�����nh�9:=&�M �|7P�q�����? �MW��������L[��n/`�RGd�����ٿ��Km&!�e�V�ʷ��eS��\|��O��_�k��K�-5�y�g^ΎIoo�/�`,@��s+[7Y�/:g�*%4,�Ip��bp�1R""�����X��	G��ޥ1������Dk=,{%��#σ���GFFT+�T�����k�בG�Ʈ�:�p�`�y���
���G� `�V}�	؊3�c��%p�%�؉~������C���`���Q���!a�����ǥ�|�ǅpcW�V|�tڡ�p�mm���2�o##q�/�y�xC��(P�*���S]����/��I�)l�:��6�zW�6�uMa׋uhD'� ���͌]��N�dk�k�Q� ���T���h�Iܾ�a'�%~xS&c�1�? ��s���HԻ�y���	a�����"1e���F�g-6]���t�)�Y��6�(�c|��+��h��?c{LT��`S��y�ߴ9���"���������
�F�LMK�͂�?��d"r|\��AEM�O�cۭ ۇE�c�G��_�,Fe� ��'�+�����*��G�B{��'�Οq$4��Z�-���֒�x�R6{�
�u��;)l7)�y(���8���fbB�����0ls0h���a���֟�V�����w��ڢ^�����A�'��ح/���DD(�ِ]=TYi*���<1�O���P�z�����ƥ�٫*�0ޢ3J<4�Z��B|`�4�"�_+���chc�b����Vĕ�RV�ы춐7���R�I=�Q�.U�JK�a 'z���9�_������F�{��>/��6�θCu���K�*�ϲ�n�������@�_������^�Tܡ��˞8�5��ż�Ͷ!ׄ B�<:9�]�c��2��~H�p��`�u�=�I�I{� �	F$��:���*�����η��^yt�R���	1}�L9@Vz׾�Ԩ~ͧR��u�K��O7�33���&'��[�up0�Hh�J�7�͇L�Q��Q��D����)9;�GEr;�t~z�l�y΂D
��c��H������	i)ߐ��Ր�eȖ��J$J��d2���h��q�y��)�J�-kvIw�W�E"�K+y�=Dʂ�y_���kkkW6�{}p�O]]%�>{��E��Lb�5�|$�����fws�I����I��ʷ,��"C\A7��h���Λ�ՠ��d�	���t�J�J�:�p�ܟmǡl[��Fѫ�  
��㹺��l�h�"���gJ5�l �f�A���2�#֛.�eY��Y���B/��v�N�Qqи���c�G�?�����Z8��ẚ��l� [>'t2P#G9�0l�!�����4y@�
D��[:E�
g�ps�EO.����skR8���^�d֘t�S���Pd$�[�60GE 4�S)��+qe�x�86_1�u������f�m�HV��V=iՑI��y�����������Oyt���_-HVP)kx�j��ũ,6\d��&OE�z���Cg��~3�{���ME�
���m�c���ۛ� Gh�S���qwm&��W��t)'U��3%�	t��1�o�ߍ8�~��ճ��x�uU�Ŧ�g��r忭U:��hii����=��&��7a�l�Ȩ��*���~ =�9�w۫�
��Կ��-�WP[k��$�����jL���P�lS�P����1��ah���w<����Z�Ӿݮ�S#�k�4�7)�K�C����l���V�Ѵ�b�=����7]��e�'��<����*'�\l'�(ˢ�o�Hp��=��"�`MbM�bӊ�죖�|���pb,�s��;3N����C��-X��ggI5nW�������A�>��ec��/�L����~gT7ח�h\ �YI�l�L�d)s�p0Cx����#z}B���׳I�j���	p�ˣ��,�Y:���f�&4k!~~�h�蔁B5¬�0�����]=jlǴ� ��o �������%���+uU����k�����;++M5�,A�W�~���L�4��?:����r;|Sz��βl�}���`lΑ�/v�����`� @ÏR5㽱M���칛���Y~=XY��"�`�I��{������V.���#i��+�\��a��5'.�'����O�~�eG=�z���b��;Y>ĬJ���>-����Bkg�|���/c�>��7�iW	U})���A�>݁�QӃ����[.�I�v�(=����Q�#����,-_'�([(�JK�,�(0���6K�s2���>[��Gs�B��_P�JKI�}�D�иk��gVFhf5��bcf���vC8;�դ&',[���&ly��	��:U�:biQ�q�a��Sv��>�L˞\p}�8(433���e�7)#�V��mo)'��0�m���v�G�ι�9���2Y������(����>�d�� *���1	e��uus�@�ZO���es�MOT�`Ѻq-��'���%*�b{��HB7�H�o��;�#	�S�[YZ�.M�NOei7�g�����m���ʌ����m��d�.M���<�M��m>�MbUL��S����=#��o�$��� #
��b2*/�����).��R:��v�������pi����jGǜ�d��~��9�{w⾵���x8�{��c�
�y�iRTem��xG3��ݩP�b���G�O�K��|�w��+���:�:}tH��P���P�y���q�\n *L�h��{��ƿN��8M�ƭ��q0/�_�V�u�ѻR�
��/e�ў����V�,6�UexǨ�`�R�L��@2�zZo�,-������F�Rp ��><S
�4�D��t�����L��ك`z{{K�ʔ��2�W�eXi
'��<#)V�H�"�2 �{�a����y�У0�)�SS�eƯ�us����8���x�`���*eF�7h<]�����tH���@[��ZZ������6���9��`��VT`;!�[3I������3�@r�l]��)g�J[�%	���C�g�t�g�RR˅�� �&Q���;ʯٚ⡞ț��M_���Ey=������U����i]@�M���	�#F��gA)@|d����d�M!�C��#}�_ˏ�t}���dgAM�A]�<�-�8===e�=��Ѣ�U1���k#����?>@L@!�~h����6���F[ӆX}NZe}N���(װ`a	�N󔚝x��4�#����$�;���`���Ll�W��%"$��
i���2���uSf��������C����\o���ņ�0`خ�{�ɢ�ַ�#?7�S8�?ց(��VyD��9��ђ�>���b���W2Q��.Z�ܲ�ۖ)�	�k���L4l��*���J��y����Ɋ�,��ja�H���
�y��hr�
ǟ��=w����qL����R�!�c�wUg��Y���:^`}1����
S�	�V�P����#�b�o��>��N�����CL���]^ma0��NƮ�g��6-o�k8!$�?����0�k��(��E�ީT�rg>��]EPlk���ZAq���|	��6>{������X�j:�84vxF��:�ۢQ���G6�V��V��U�f��8�ɡ��!�ɝ-B��#�PsPl�����G���m����5&�f;��)"��(L�Nk��`<4�:E4sA޺q�1�E��66tu����tڮ:�d-5&"�lM�$;0ת�}���\c~�J�n�%�'�N᳛1��6��{���k��K�|�S��u-�T�_���-l��� ��p9[�p��ॆ.�l��WY��<�y|����@��Jf�?�n������:^]25������e��;\�������_�t��^Be)x_�w/N����w�$��q��<%����7�ʗ�]��2G�j�(�>�.d�<��w�V"v��t{&�폭jC�����'x�s�+�Y�_����Ip�Sw�9@�3j��}�x�@��#��~��/ǅF3�b�����~����\���@����̄�%)WfG�ș\+E���cr!H.��`�Q�����S[����x�l��h� ��5D�ඊE#�_
+
��T���֯_j�z����d�(n*���C�&�g]c�j���}����Z�])%ɍw�	s�b̙r�9r"����C:P���u�@�d>�=^-�?��@\<��_f���+k6���E�C킁�����鹾����(�7�����.��<����C�����'6 ����	��]z��TB&:릅_�q��a廉���^lU᧬�9��'vP9r�������`c]�k�0u42;S9y��\�{C闫V��ƮG�M�Asrh�[D�$�� �)��| .�~BZ�8��+"BITi�q�ɳ�e��^���p8�(͢m	��Y�N�����^L�_�N��lk�&��qے0=�/��cX-l<[���Ur��償f�aYĔl�|��\��l��OþU.x�a<:1��%ø�߬o��3��X�E�,���l��=�-֡?��c����v�FO�6�M4z�u7�W�TB���䤯}r��Z��G�O�n�
'_>A�{��Z�u����Ä�ٶ �gur�_�ڮ'�|�y�3ٙSV�������ț�����ڷ����GLR3v�~1�0�\ԯi1t��u����GT��-�_��+��c���">*G1�8����H����y:�G������M�FM]��a�Q^�2��壯�8���֯?���?�y�z8�F��e?���9摊o5L@-	�(�z&m13P#n�߀w3��������jh;_��J+����.���r	���fq�+Cg����ͣ�����mJx���.jG��&���QI�rտ˞ �p'�G1�/QI���������홺<4�{¹�U"Q�sw��wm��\��,�R�ƫE9#�o���ߚ�=P�S�˵P��(i��]��f��qIn���Ee�Zz�좒F��̌�q�T��P[�|��<���[�+�pu�EB�	��!l��|�H4>X��ۍ 3Ɔ��z���U�m欼��D��l�h� �>8ĝ��u��q�hc����VB����z�WG�YX�/]���@�Z�s|ѐd��-�BE뮤�}2i�J�SH��%Ҳ�@ ÿ?!"��23#N7�m8�2�2Ha��ne��Z�����Ӻ�C'��D�v�� t�s��t3�����t��Je�6˵��L�	$�u
��J���_����^썀��V-2�W���h��Cknnm����`~a��T�+e��OB��?ңL^����w�u#yS�ы��[_��������.X%ʤ�]�AeZ��y���l,hiaj� Rn�SL�d��|�e#��|��X%����y۠ �I&�?�r?|e��> � [�>�!d��ө�!�ꎃ��j�s���I?YV�
�p"	�������(���$p9����� gM�������Z|�8��	�߬�^_�@-�o�<���������Fq9�=*h jz�@`���}u531/���s������zR#AOXɉ���p��q�]"�+C]\n���zX�/��7)lk�h�N��-��=�@���o���ۍ�����$�i1$��2P�����TP	�%;8��'��QN?d��'$4�K���UO1;'n)��[�y��90����U�b� �X�Il,�������2Vë~b���9.t����Tdh =��i>�uM�"X�f���b��>,^�j^�E�V\Rb'�`����w=-}^g'{��R�~�̩�́Y���sP��=��zII5��}�'���%P?��+C�ݥ12����ʈM�ݐ�?,�o��f�h�<R�T�/�x����w4W�ZgR��?2�̬ʏ�Bo��}���( �կD���w�&�.�% d�n@�����=�2H0���,&�%r���B���x|uu���X9���74`��������\�jB����Vj=}�L�.�Q��}Kӗ�^�˪����]B�����S�$�(��U[��&����n6i,^v�Bf�)`2ޣ!�����Y�mw������D��?xx�DYb�<M'%Cΰ��L��@)w���ѵ5M��?��?�w�'���\gw�?J�[�%!���s�/q~ M~u	?��?�N���i;5����R�@�D�bߔی��~U ���@������^	�Y���{�>/������^yt�n8+[��q��naB���W� �����w�}44g$0þ ����e�"tF��S-��GS����D�1�o�vV�rY:�'ɍc�ʴ�S�����6�w���z��0l���3AA���r����ԉ�7ס�3όʖڂ�s� �KA�Fu�������;�%��9g�����>�B��9��v�U���v�o�$,+s��oc N0s�I7�4�z��n�w���u������W���Wy��D�p~�+�|B���iǃ��OTt�V�����{���M\s۔=������Nb����Cr��e��������R�U�����v���;�wy���rk������R1א��صq���,��G@ٷeD`�m6���)�`k�ut��f?�B{���
��mftr2&-m��B�4&�;�h�:$CS��mZ}��x�?�á˃7-$P*��)��'�L�!Y��ո��v�(k�Ŗ$��E�!R�AF��$�F���tMas��|�z������FAj�S��$�z38�'�� �{4�>���Y'�\i~l\���^�"�_�#o���bs�Y��o�8)��?�W�&!�x>�#��(���`�O�$N�W����W��+��*����w�e�����N�%��k� ���1�ݟ�ރ�S��W��P��f~��<���w�z_�-h+�4j����_סW��r�ˋ��x҆�5�B`z��>W`�p_��������ի��V,ua`b���KsKV��Ak�L��!���z>�;����^����GU��PMQ!�C�vE-�Ul���+���.��X��=�=����nb���*�;ZwMOLD�ȷ��Ԭ�ac�99�&՘cX�@7�����R��b;77���I����-'��¶-o���;X��m�M
��y��?qv�F)����EʪWK���JV�
�XqSK�����{�%l�5==��qi;�&�
��}����X ��C���rppk����2��.��G++M��X'ց�S��/a��P��p;l+��;��f�3KK�� l�6�iC||�Go�jv����v�Y�{"磋��N9r	��=O�$ w�Bb<ܫ���=q�k��g # ��l������7���m�z��;�8j�|��yL�������R�!բ`e���M���4�uXQuw���g�pc	c��'5��9�b�C�����n�W<�F�ɧ��7����ݬ���b-"qt�����>~�n:�M7G!q!`��{�WS�������>���`/kE>n#"(��#�1{W=4�=�����}�z)�����R�P:*DӃr��([L
{�M��ggG.#�����2�sX�[����o��TI1�R8)8�Y�:bhD�]EY���#a�`ūRwlF�.�8��\�N]@�[d娓���sli����t.�03�����D�[�drC�^��2KNM��}��'S � �	;��ɋJL2��M��M�?�ؕ�����hV��h���zZ>=�JR�>��3�3�U�+�"C���g�RN�e���!�=���9�;;��W�Hh��%�?��O���M	oq+�����N0���vISv�ޡu�I�|������>F�,�2*?cS��Hb��rÂ��ؔ+�n,�$A�E��G���?;F���sJOJ+�S�(��@e)J��f�3[	ޱ��tܽB�\#L�4ǳ,�Rؒy�C/�����'k��[o߽[��X�\�Mi���;�r�KԁɆ�t�J0�N}7�Ɲ<�j8�x���Q �ூ���G����0s�.�Ud�Vi?�Gi�e9���^��Uʺc�q�&WL��*�}�[xk�-��J�����)�����v%�je~����������:E�MM���
'\B.����!wI8! r���a���P���lݺ�:�U�GE}qG����٤܇@{��֢��ńfW���W�?#v�)���-,�-g�\!΀�=�P;�oH�	ƿ��ȱ�.#&QҪ�X��j�2UK��rd�[8p�"��nM�y߻J+B�!�3�ӹ58��G%u�E%$�2?�G匍��iW3� !�2cҲg4��x�<�L�vyc�Je�*����ﱁ8��2c�>��A�9�3��vV��o��D���=�Q`W0���٬��u����i?�:�'^������!�B�HZ66�
���� �t)5E,u���3G��V/!�7�Ux���%����`��|F��UA������x?Ȩl����Ms���3���8�ť�R���1bb$��F�?����,i�=|�FO�۲ $�ƄOah�����8��/&�.Lj\�j\��b4���=g����׊ܑ<�$�>JXT)�_O�\6�W��'>�v^EvT��ՠj=�C��*%��}�Pt��&�+��(�k���!(�3lw���ب�b%��;��TV=�l�D��6yl��l]�C@�m��5�d�b�VVO���ň|7���y�O�f��6�l������a
�Pq�}R�Us�`������]6��<=9������I�����"�<k�V����r~����<���|��
}d��`m�iw��t�U�C�������H?��" ҷ1�g��!&�$q��fuSućy���_9E�y555����.	���v�'�c*\�TO��Û�[���5�)�"S����*�~z�ewf�M����2ju�X���!	��Uճh�r�y�'cN��/����0�#͉��֙��Ъ�W/��Վ(�(��:�[D��ﯕQ������Yc�*wa#� 	�l�ɩ)�ǁ٣���Eo��^P�=*�e��>��wg������,_�N*�7�B>a�'������3�ƪc���ި�vRp��� �zm�<Z�p�QL�G���x��U,T����B�t����P+�����$��̔��sS��B1��|:�/����W���8]�1���uYN��Em����l�fX��@s�9��.ew~�.�4�w���c��5�5��?o�~��
7���I^�ޱ��sXZ��=;��RW�4�i���k�<m���q�a�~�	�3O�@�� ڏk�o܅dU�.�i�ou	�ǲ���$gA�C�֥ҏ�*O�r"�6�$_]��~i�mY�C:U��ߟ.�����)��7ǌSV��ӝ��^�����"��˩�SkT���ɹ����n�p�~���	1���ݗ ����}+GZ�ؼ�ߠ��P6�o���{[��׾���JEc�M�[7v�W�[S����ν�(�H��E���ܛ�\�p�_o� -V������ev��tDFi;��ǌ ��"*�~	���F>�G�.Q�f�	�}	�U�$�����.�C�p�ax������~ F�턆mm��ym���e��X|l�:�%2b%��l,�M5s�f����e�u٪�@Ӓ��ު��M�b.G�ґ[O�(M��$L���Vs�yBj�����6g���B�dkG�<D��lkm3�Q�g3KK�2�<�lU�-�g��a@���t�1��ata���TD(0ϘOyxy�[�����B� ��*o�1q�ʙM��S�f�uՖ���T�����o�L������31WiK���?�P��[f��W�>�cD��Ϟ�Yj���sgmѳ�������Y^� X���{�u��E��
�H֡��Nb�㯄� -����=}�VI�1���͝��t��:��1��1�?���kpO9�����j/Ln_+�w�R*
�V|�T��[���N�cD�y���Ao��d9	�m�����QЭ�tuu}E*%�,E� 9�`�F�c��g1* צjO���*����6�Q��h��D~�.ptr�t\8��y}<1���~�CSW�^���V5^+nQr�:���U��#�k��&��.����(��?^���J7w�￴K��c��+

�K���FΗ�ßZ�a7+�p����N� M˷'��S�	�J����5;�~��	��r_�]'�`	�/��Y��_.��E0����TO	�Җ�|4۸+����Q�l'��.^�_����Y�EE|�tu�d��?uQ�7��1��]i:XWh䱡�%�4��2����z�WD�-�ΘbP��E ts�����5�� t�+�&zu�?����߿����O��cY~!!577Al�TKe{�� Clz��R�&�.H���R%M��g���9a��8�)+��<U�����F> �X�;������_�0��K>��|���,\J���ݪ?��UY���w[-�_�qE���>��}-<�hTfbb���i;	_.���1c�@�57C��U.||B���6�訡f���S:c�2������o-�����C	�qa�������?���Ur��b��K�����[<�w~'YH��3%EGni���;|u�)����J'M�BC�d��$74H	��[�|���Wl����;R-�m�*��c�D�\��0��{�A�1J�.�,��@����^�{��4�,��rb<z����ҵO
X;���G9�2�1�R�諆}pL��+�C��ʭ�;ޡ��&
>u ]Њ^����J>>�Hi�fq��r�� s�����ђ�D���ؤ�C4� ytu��'��J�|	���h;o:Av��e�$��M/�U���D��E��ig��jۋ�����Z�љ�j~Z�$��B�K�bg��#�WA����Cp�M�=�A�/b��݀Fdp�y�`�%�����,A���9�`����In%���넄̴w������B����� ��><)t6v-j
��Z�-�=����2�k)E˳���s����.,�Q�
w�wP7��#��Ps�h"vn\K�eo����+��W.��q>t�����ۺ���.~�>��[�I��� :���J@�1�ʃ7�ŝx�f���C�_$���L��[�|'���csQ�>��kjjz_�$ommE<�ka@ ���Q�
մ(3�p�)//��w��~v�^�?��a[Og��/c�>?�f�f{`k'Q�g��۾�~�"zd�l`���ެ� �9:��h�g8�o�m�2�6}��\��ƯtA��~a��o'���5�+A̬��x�̷1c�����~9/��+���<G�4H�Y8e2(:9�����@e-݋�U�;��"���<��	��K�������k��}�Uf���H��}W�H�+U=�5`g�;���Ÿ��k�&���K�&M����9���p���>�.���� Ħ�F ��r�B�����{��A��O�<�ՠ��u�C������&I�t�lw~�O:9���#v�#^��9�2���F��o D��mW1��	/�k����X���ra&�Aew�Ư�\�F��x��.��؉.���q��PY��#
7��R���ȣ�u������b|ͮb��ѹ���T�N�b�&�JU���p60�e���Ǵ������/�����ɱ�
�>�)�l�h�Cw!�wCocm�v�4x{��(��= \����G�^��O���gcZ ��cJ	���R	ۈ�p
����bT�x�.̡`�����X���L��F�f�����sG��5y�Uvް>~�x(��}O��E��7!�L#H�+E�7���)�8�Ƥ��XQN��s�A�ORx4��Hm�㫭��#��MM��~�l_�O����Ԗ�����	[;�ck�ž���MOwXh�`�����Klmo���G*^����g�1��Z�����*ᠱE��m�
��*K�� �04<L�b�C��`����4���<,���c]C�90Si��'��`g`�R��}���s	Q�D��wk�#�=�-�E:�J�"��B�� ��>/����K S!�{��m@��"�K��3E<l<++ˠ|l=ӹYG��j�PD��zJ稐����N"m�j�I[����Ѭa<- @Y@Ц���[آ4�����ݱd�v��k|��)˳�<1�Ҕ�ӕV8b�>�SP���T�8X��L�J�m��'E�����G>m�urv~�aX6vã���tD�*��t��)�6���S/�X9%��1��J"͎�pa��^i��Չ���%��l�p6՞��@//v�>��5u.{�!�=^�5�ٱ�#��s�����&�RJCS��_a����?]�U#[{�2.ט�Nv�b�=Q)7����e�X�g�F�������'�E��n.��0A�^�{o{C�K����p�+u�@LQ�7*l���,!FNm����Ȫ����D���'\���j���4�� ��Ii�oߖ}�.�~��XQ���k�IcYOS|��G6���ׂ����|sl����{jA6�3�sd�!r��|��d�r���ٸ�ō>�I��QE|��eL�!�0�-�~/�o� M\y�`� 'V5
���n���e �4��~�z�=����:�;h�y�!z�+��{N������ �w9+���{CO��e`@���O?����b�1/��>8x�Ն=s>o(��w	�7�˭q�}�����(i��	�};t��
з��f�2+N�+&��}�,��O��bk�>E�_���*���>�Ƚ���z'qH��|���tk%� iC���8����~eZ��ʉM%{ǖ`� �%��J`!~��	d4��۬|"�{P�zQ����Ӫ���)�~	|r�芙S&ʠ�$S�y�ޛ �9�15���ٟR�8վ'!���fH�B�z���tɊq�%������	�O�^�[��/�S}jl���А,����U�*��X�V\O��ց�i���k��q���y�}0
�Ʒk��֦����wc]J�!����@xa�R��o�+!ٺ=��*Eƾ�'MK��u+��B��=Yڒr��n�YW�  k��?SU��N(��-l;u����ǘЦϞ�����u�!R�����f���O�J�J`z�m�y�6bӘ��f>��w�fk ��l�A��5����h�b�kr�� �#��$GPZUN�8L��ͣ�'lh����C-�Woe���t��4H�tJ�t�4��� 14�H�t��C���������9����O����k��<k���i+��������9Q�1_�>��[(*�떳������}�  ��עk���B�7�����c.��/'=���Ge���[Z~ �G�X\N,���jF�������4�?}2��;ZՌ�
3������1�R6�xI�(*T�'��O~T�,� l)`q������I�������%��ܓR��y~�p\�-���gN��T�>�(��
�W���DC��;��C��%D�70P֍�9H{���~�Le<���:�"�����B��;�4V,̽���U+ai��E�����?�\U~�l�f#W���bN�\�g`���q�%v�"�IUX/zX��iO�oRo�
C���o���Y�.)���f�X[��/��=~���@d����AA2� 󈈋r� �V�E|��GM�$����W�R>���p�CO���d{���*�α� [�N�g��y�kg���nP����H�9�/�\#33����w���k^�+�F2 ���33�b�o��dO�y�G��=��ZF5�`��_�b�[�����yM�MV�"CM8+|����w�V�6O:*"]�ƚ�AY.2"�R�h4�ԕ��i�v���1O8%M����_���S�$X�;��ww�bãAM
ņ]�1� SI�0��ܓ�i�R�P�$�N�9�6���5E��<���*�2�-roL�٥s|���ӴXf�!�v�l@uOi8�́_a8SC�7���s���4��/?n��k�����'`7T���+))9�e�����f]ť���L�k�yX�Knю�wh{w�Ш�VVC�:�ϯGV�n����JI�%�'�p`����ht��ٻ?;9��r>������ mI�?�����'�8>~2���`����)W;QQcד�3��i?0�����E�����&z�+��&�6�N��:���6������t!�MB��o�2��FX�h	��m�8��P�i蘔��e�(���]͖�"�x$؆�m}��L���t�^`�$Dvs>@S���h*]�?.�J1WQ11��I���
7��ĥKX߾�V}�dC�[i�;�&$�U�L��	9�`����{,��j����%��MD?�����V��+�4-�74dT[� �y�4骪ҶrJ��
F/�ˣ�!قU���PbG��KKK�I2�m��Vξ���}���R @��g�Ss���6��ߖ��u^X"�����n�8M#�2KZ�����+������2�-�{��o�!&�k=�׹�*S����M:\_mB��WN�C�*�Y���!�/�]kG��Y���0��9�<� ԡ�I4	a�b����N�6�2�Y:^��_�$�CҢG H����������m��d�I�0�Z�g��D�Y&U��2�i�U���D(��(�9��v
v�����N��t��6p���`���I��v���� �z4x����?*׌���|��\dG:������a(XX����W
BC�X?=g9��
����*SC��l�Ү��g1��i�	8�����*��47`��%���9P�I��0y�".Z8=����zq�Vݤ�J�y�#���^h������~�1B�?��X�x5B���'@&lWTL<`A��Z[{��+٥VEu������������`�t�{���䚊K�k��u��7�E����W��F���N܃�^��
����]���🞟6��0Ƅoo�9fO �p���:�@s��h�ZYX�R���3���tZ��d(HT9�Q��uʳ⑱����;�UP�6]��b�)O�;��ܶO}��'y��Bk��]��XO/i���jDn�UY�p�n隬�t<@M��/v,8��v2�H&���^���^��Rs{}����_�i`��D�ܽلػK�89xI��)3ͯxq�V����~��O-C[��X��*xzd��n#n��M�]?#X��G��c��Y%7~&=����y��0����_)���}�o��&�����z0��H~�8�2�}�+Gf!�9$}>��Dzs��F~�/`���Wѻ*qe��̈�#�U�-�p����|\�C��j_4�R�2A�ǂM�-����~�0-�DF��R�!�Mo����������s����;���ܜ}͟:I#zNl�n��@�`��tG �ʘ'<�,���e�������[ m����+pw��u>���n�bj������D6�r ��.�
v�C���q�?+(��=��:�?=�� �E�'US6��� U��F�?�j���޹���K|�f<��#CK�r�gnq�̨|�̞C��^������*�\t^���o�dl�Ua�A;j��--��֢������'��V�۞�E��ߡ���̕F��=ѓޓrjj�,ۡ�6/��������r�Y�m���m�G��҇��~�'���WN����ϕe�B9����;*']O����;hy��HL&'!~����&&xĤ��?���旓 5���l�0����X.~�h�b*�����UmZ��<>���{�+0���%u��L}aV����'Q�
�쒑OZ��
z�E:ڋ����>z|�V�E��-�CL��@OڳwFح��,xª�����
���قU�BI���O4��ڞE�,ȝ���W|բ�ۈ��AU�K���@"�X�_�#��B�dѫM\���6�g�$���F��W@f�x�<Ȱ��Ӑ���&��4ʥ�s�2+�
��_�4��nb��(1��?�W�F%�2�b��E�H�MyBCH�1���/,��Ɋ�MP���t$$"zL���4�Y�ء���I�`>���(����(��%��E�:�,�uAGy�+ B��;�E��E�|}ܧ�$�LA�KYM�K>M�l��&��l|��g���K����lix�$g�O����m#�H5����ș4����:ĿTd��鯸��)>��
<oXm��S5[���ڪ�"`��>D��BLcy���J��ot��ED`~���~K	�U�^�"�4�B�w_�l��I@w5�V!am���G��y��a��H��1M(Ҫŏ�WDۋ�;jY�����I�=��z�$~y�z�-eU_�6ob^ErG��Br�5���C?��^	?Z�;.����-��m���E%��e�>Yd�3�b"��v��8 sK��6|xF�mShp64����:;?����eV���wE}� \�-��~W𬯯��cj�v^���J3|����K	;�y��2�d*g ���Z_������ϯm[�({�<�/�z�1���� K,�|VHn�-���4�n��JUӅ;�Xf�H�cg�$ q�q+	��#�W��M5֕"dR|6ۉ�)+�faǱ�GkI���KKq$<�0k��3�}�t�B�z���-�%X4Q���889u9wʺ�qQ���\&���؇� ��y�s�S�ӑB�3|	?�W� ��B]#q�)��+�?�"�é�/N5���}�+2L�z�1�u6r�|M�=c6S]U���2�N�4�[6��y�4���tw=���f93�F$�à�fph�uZ��˞���I%�A�P��9�=p+ŷH�&�^8�먳��e��-5GO廓0��v�)|��,#�4%2!�;J��穄D���r�M�m���$@j���[n����`G��S������ގζ�˷ ���|�����Z�EJW�U���wG���:,N�cy�������>��q� @���=�ef��!�<c����D��ʈ�f���57��;hTٮU�ش0�"�UkN�Ȃ�6���D�(���2�&U�/'�B�<mM:7!�?w	���׻"��9oP���|B�W�Ю͈�'X��%`80��-Mv�nrr0����N<�\W���V�5�6���ZyK؇���,h��J�y��䵵�Н��1�I�!i�1�^2)�<[>tu.���]o=@T�ى����ȇC�(@y#]�hRSr�f�8B��k8�.;�u!��BƵ��~%�I�q���R;+JJ�ל&ǆ�y�@��(�$S���GZ�FR�>�[	�r&�U�|�a���fM�����Ϛ�FV7`EEE�9�-�*�0�k�-��H��y��/%��}��E�[>~���߯�ʓn��;��Z�^A�����W�����R(8�r��nz�<���1�"��4�аL�Ԥ{��Z�ue��������z�#5Uc�gR(�8��W���h;^2d<�
�.���M��*L"]�9\U��F�:��MM3�P�����㑐q
7�j����	T7�}͚��H����S&t3I��9#`T<<��{���΢q�2��E5j��۪��Zwr��[MɊ���(Y'�B���;";H`_ೋ�7���9}wZ����~�h����;��n;K� �n�.�R������u��n��@n[����tU1>�G��hgggtb�-1�`%8U+��֞e�A�y��=J`Qr�m)=�m��5L�A��'$���zw,m�Z�R�!�X�F�5�i�ט0%�L\cU��:�5�/�of8x/tYAHh���i�scc%�/�s��Ih� Z�a�X�f�h{N;2���EAO��5�o�T�54M�蛩4�19^Y\��,��l��qƄ<	��B�_b��O���c���绻n�b���Dx����˜�ƜJJ�Sn�B.�>%cn{$ёk|^u�`��?)Bll�7W�'�s���j�e�\�優�0�b��O2���7x���3 ��r�n��cS>��an;�?j�Z,��R9��S���8������p��f�Dd�\z�T�̫�lrwQ9ܔZ��Jt;�L��<�V ��F��@ ���&�����~/�6�@�y{M�{�t��4f+��Na����cH=�"�o7�FEQ�"�XX ����j��� �d��#MO��P�k^F����K,��8�NF@q��t?�\��4��D�*�y���,q0���lG
Qٖ*���P���!={��Z�y�U�Ņ��5������KR�a<�S`Am��д4�j��޼ �b=�r�yu���J}��1Ԅ	����g4�ʋ���]�����v�'��p�h��}�*ħ �k�I�m����E ;��TA�t�����صz����'*&��+�����G��ם��w	b4T�s��߷�9���<M�b~�9N���[+}��cx0�*u�#��{�fGAM������bZ[��}_eX?Wu�}qd��Sn�"L-JE6��i8�igL��"������R�19�tmW��]&1,'M�E�}��z�+��d����+�c;)����e4] le5�a`����6=sS�Iv�)ߴ2_��4�GŽ}���F�����:f��簔PMb��,����麠a�-wt��|��	��UTO�_�Fj�A��e8z9��Ap�x��)S\\ܾEq�y5+=q�����@�q�˷��N׺�����8$d�o���ꊊ,E��1X-չ�R��f���Y��X���>!��S��N�z��U87��bc��P�XNv6)!&&	(�� ��t�0����=�\lί�76���L��R/��j8c�w+�@����ts��ˏ䶁}�����^rkii�BA�6(�Kd�,��Q緓����ؽ�i��;�?�W��Z�q-z/�h�^����_��s�'hl�����6��:�&�S�)��	� yit4"6�;� �>f�=���F*�b�(�	I�������)q��~���ʣ�����B�O�T|�f(�rb&���5�8�STR*#(A�}��@1����嵟ㆬ�_�x%%��c>G�J����1��x��v��@C�1¼�� ��0?�2+&<� �\w�j�
<x4{�c9�=�!�����𳚵�]���U�}���;�x�kmCÛ�`W|�I���ً�з��~,�_��&m���꺸�lnn�d�4UEE��x���e�h�A�iauun��#��W�B�<c��<j^�*���<�Խ��-��ZoA~2��bT���H'c'���p"��ډB=(HκʬN	\t��&���ss�(I���N�����	�-
�o�d����xVc���MdQ$�:��ֹ���#8)��.���V|��LL1���UTH�`���1�t�`Ĩ�d�j������R2��Qa�PX�����Mx& �fη�17���=����<�z14�a�� 3���9��M��5��-H�O�\���
C����� �}xR�k����[�_l���_���m�_�����l<.�vpu�:ߏ�t,��I���&���Arr���;6��W��x����s��X�Z�o���5D�jA-��fu���S##n�Nil^��s�X����"<<�Bk�_i|6q�ڙ>�+zY���m*�������Ufx0%�.�t�h3Q-w��z���MM�z��э�F��U��m������K�4�D��� ���9���S��_�l�vڷn�	 H��Yd�ũ�]�6�=�����J��R����t]���K��E<*&iK���S�ݞ��3����*L��Ӌ���(4����P*7�Un
�k�'��o=���n�WLdg��&�P����ZUx(u||���y��(�(��|���E��JcC���J��Ī�^t�nfH��S�0���}�å�n��+�a�;�NMV����#sKj&�u..���Cə�o-.��so�X�6-k���!,hj�^������	��9I�v���������::Ў�\���ϱ�M�{I2���LL�g�?��.��1�,�7�>+VT����r���9 �����*�`���f.z�F� �~s,*&^PS�'ۤ1�#N O|0x�s�o������by������4�xl
�͹cS'����ٔ�߹s����㕵�NY��Ȃ�
 R[<�e����׃����k��r���hc,:���p~��b6�j��u�t;d���
��W(��F�&Am��Ԭ�A?��|�M�R��ə_S�OO���啕]9K��"""}CC���@�������t�Le��͕�\U��Ի�t|T�q0�6(DŪ��'�<�v}���(�?�I��hZG����l}�N�D�a9�g���95�"gȑ��Z1[0zԁ�bm�
 n��' �����,�N�A��巆�o'_FX
�(囡Z|M��$�?��		i��u��f���������;+b���0)6����I.O.�V�`Q�U;{�Z`�'�_�~`��\+/��O6y����'���l�l�>������R�\l��χ#�Q0M�:'�B[�fӇ憳��v�F*��x��Dz/bȱ{@���fZ�3Ղ���0���4++K���v~�Se�֋zG"ӚP��0��뱈�y[��>���S΋��t1�w��z>m�4�e���J
�nogJOO_L�$b��;�|����47�2���x���!O���kiM��]��E��ˠ'�%�H�)Y�d)$Y+�ʆE�����[ۛ��z����a�Yg[y�Eӝ����mȟ�ү Ne0�0l~O�����T��`�***G� ²��� @��|���,�_{{*Xt2�>AaaL<����%'Ei�q^$���Z2#����^��6��u��II.�&=$*̥�aC�����U����|�ޕ����`X~\DD�@�ދ��5R߬�ʙ[�j��5ς(�:��?�b�}��i���0u߂Q�}B�Z�e�\�ss<暜�WWן']a{�lo�s�a]�7O������ڽװ���c6K�-�D�r�~B�֕ssʥ#Z[[魬���EH�F�o!T-��˒C� M5�g%�r/�`C�Ws?��8�i|��gʰ�mkG"PdK��Z��U���R��4�3(�$A����.���M^���
���`�xM���ׯ#l��6���|�[�9}oB��]���bs��^sd
�y��l�#h�It�w���eE�G����G5qLT����Q���9K���o�l1���}`^;���b"��i���+7Y"[[B�i�Đ]MO7�_��ʘ�� Oe֔�E����6�T��e��E��|k�o�fe��\��e��B�^�~kx���g>C�6[�k�����d�kͻ3�����봧�:2���?�U�w7rv�P3��L�=�,�f�hWqC94u�ώԙ�_|���,��7��Ԛ�J� �JZn)��hq�� �}����d���������𵮤��ZŨ����kT����l|�B���5cI&Z��eD�iK�+��4��LC��a�<Rɶ���a�G�t�Q_$[*���(.aK"�2����S��1~q���_� T�oX۵ �H���L˥ruONO���,,,�t�Q#��@m�ɺ����l?�e���b��(��|���^����6��$6��Fig 3MG�@���/cTe��Be�흩*JYB��X���8����ϟ��08��5���'^�����_�#L��^�����:S����Y�����Snnt���R�S�k�D��uud~2�71�P�Nq�mBH�"J9
��~9Dt�3'�T�
T�ɟ�v=�y���cbb�B��Ռj뒡�A?^O����j4���:{']슨kƤޣkD^��`_�'kJ����(����I�G�j�0�k�# ^cӞx�ߞ���D�
ٺ�ִ�I������P"�/��R�o�ovq�Z��3TA�Ɍ	jGg��T�:�EX�����
	GN�s@�����[潶�؁17��ԙi_���|�ї�V�\nx8���>n��@��'�a՟�r�)�qUZ	%��M-1ʠ ��}p=iSs�m�95��6����/o.���n���{��h�!x�������C��R�$1��g�(�884����8�c��m���o�}��!�5΢xK��P�ͭ�wwvqa������0���������+�s�<��Rb>���o��8�����\l:�����xf�ߘ���A�QmKGK����oi�^���z���4�ꍊ	1�l���q����q:/.�z��4���lR�EE����؆/����.=c���;:�<4��	�2�<=��0�@��y,��<�a(���ڍT2��/��%�6���~j�������)f�&,�V���J}�A%�69-�*��?�w��PUzt]�Ͱb"��m7�D_�< ��$��Z)�h���ٜ��7L���D+@F$��x|�a�Ս5�	��yY5�ݦub��~(���
��	n��o�կ}��۱s�'�������6;@j	�)��_&���+�ؐ'���22ª���EHB�:I�������γ����G��cI���f�Փ���~|�����G[��}��ANޙ�0�q-xҵ"/��#?�Ȗ��f>�����uz��v�ѝ`ZF��d������N��u�}tە��qV��H~yy&��j�o�%$,,���E�v[��}���0\AQh�a�T�r�7��ied���0��~*C���z.'r#~�������(4@۾4�6��Z�쇂V�"�K�2��-P�)T�2�?f||9�ZלXc����b�6�����hh:�,t�	���'�Çg�4�X�̉�3=�<=(8��+���Č��4�]R�`��G
���Z�]1g��T鴚�=%f�=&���;'��%$p��UL�%?��l~��
j��-����W�6E�O��_
�R��&כ��F��<��V��[8��4��v'=	"�.�}���P��R#Z�TU�ng\GD�մ��Ƅ�>���X4pXB�?n/Ot_��r�a�<�0��,��E@W]��kƕ��Q�+���5�YR���֎$��M� jw���Rަ8Ѷ��v�����0�ף��Pyro5t�́���@�Ѫ'2��t�|���&�B�i������ص?y	���7`��,�<�I6{߆O@�5!����~�x%E�׸,�Ԉ���K�F�	z���~�.�1e,FH��;ߤ�/IVW9�@���Wϋ^���<� 懲��#�T�J�h�X�eCu��@ȍ�}�ȶ�����Gd�ׯ���?x|6,�K�D
_��*?�,�Ӯi��7S�hT5 cW��H�|�����I��/"X1<s �h���)(8r��v��r�q��`_\�R�7V����FЛ����n��1�@,���"�"�4��a<�R�la�92�w�fXt-�{�d�E*�)$���!T��Cx��ۮV�k�a���=��� ��4�	|ckp�R�^;91�ʘd��F!&&�'�n.\���4:9�U��m.E=�@:\=�o#J��bf
u�R4�I	m'y�����U��V��J4M�(�켖9]��wej�bA�L�[���Y�,"+Ǻ!�H71)���JG7�zT�U�lH`��ᔇ�bn��h�He�C��Q�D��eU#�+�?�(L�()�^9)�POY�������mg�J�CHD�=���_U1)�>�D��;Z: ���fx~��xH�D�l�2&����&�_�~^C?����=9��>Rj6�T4`����Y.1�����fB'^.�j�r�% ���VVF��c��Pϋ(�!욊�0���L��¾֏>����)�i�� -�P\����
�&H���	�o�W*���u;!uH�5��8=���T݄'���Pxw���ka��f��ţ�G���}�[���k��ӣ����n��{� ���y��I���΅��i3�!t%%[�F�~���&Z+R��S�`�7����mٗr���KG��ë%��"��Ŗ�����R84��p��V�qTN ���A���Ž���v�s�(y"�&_ty��s�u���C/_�^��c�4�6�	��Y������<~�|8����ٛ$�����F�:���P65�������[d����8��W��c�*��z�S"nYL��M2�߅�rۓ��,��-�L+�L����M 4�@��s��6�#l���cI�gP�VY���~�#��w\u�70��x�X�������d/s�8|�\�i�������ө��9c�1��4H3�<�c8Fq�75؎�L�̌z�Wv���6�ieG�ˋG��v�(�vH�I�g�A�����s�����o��'�TSu)�&&(������i�:t?��o����X�c(!~xچ6~WeH��)�~���B�.�򒌌ܶ�*�X��1"����uw��%�H�p��](��bQapM�*6uG�?�n�]�~��{۫s��Zh0S-�
Y�c왘0�}+a4n���q���nA��hu�~#��m�c�х|}ܴM� Å������"z�J�5���:�4�"G��	�x#F��L�G07�'NǗF�A"����{G�d���Dv��-�A~���I_~��i�ۭr�b��3_
2�.�,f�zzޤ���"V��v~��Ua��w�|h�G1_�=�/�iQ>�9���%�9#�0����NAkZ����!�k�B������#/��G��Q��?��\iډ��l�T
_ �7��������G5��NB�� l`�� ���A趎~�����0B]ź��R0Rg�U�ۣ���&�Ӗ��`�#J=��*��G/�m�މ�MHD�(�YO'*i��`~�HD.�p�C�+���?�d������f�	�u{����W�U�r�i����*9��TW�<�,]p3Ey�,�����ue�B�}�J��C�������z�1�P�����}������5���_a�5�ٺyӻ���HO!�E�?⋇s��/�3�,�K!F\<Jv�,�s�B����ѡ䄶&���J�MX��*���}��_;۽,SM�1���M9�.��3���v�!���5`_U�:ڃ��#M\_�x���S
n��������� �ntb�M�����ұ���e��O����E}��ΊE��⛨�W593�wPG����a�cu�J����tdN2?�+B9u����We?�Q�%^�KJ���Ce�s,?������NLj��z��U+� Y�/�� �ꪘ��~{ ��?���2~ǟ#A`^	�]b�Ξ��ӝ#D���Is�9mnƴ���_��^w�!�ux>ѐ���l����ѥ%��b�L���I,�0�-�Ȭ��[�O�8M?�)���{|�z|q[�����! \�X[C�����v�(�Ă�c����6�]��Q}��cU�R���Oq�����^,qg*�b}�O�ё��|��g&<�ѯ�!O.C��H��_4^�#���īkU�&���O$2�F'��p+s���\3���D����e�.���Y��zz���_� P���M�G.�s]��P-��p&ҟ&����dV�'ŏǷ����;�Wp��{w�0�E�+�I�V,UId
͟h���W0A���-5�gk���&O�v��N)uu5!QQ6.�E0����p����iQ�G��-�1�e�j�Q,�k
L�Ճ�P���Z)�	D����a���i-��0l� jz/Zm�j�no?xF�ؐ��A񍉘���*�x��/ ���^n1m!L�Ψtܤޮ��� ��ii#΢#[�#�}�ڮ�QM�3|ߐ�/^�44��m�;>���6Ƣ��7���������V�W�^m�,�J�C¼�R4����C}S7c������i�nn�������/������B��s&��'�����%@ ������d��@d@�R���j�(p���=	%GOo~���㴿tN��婻��4!����d]����.�����7ϢP�q6r�ݩ+�4��S? L ��H��)GCC=d�����&\��_���}���^�n�[�-��vB �v�'�S.u��f�$\T�LM%wpr*�d�q|G��/O����̢��p""L�h�vT���ܡx8_�MS!5=�j�d5~˂ ���7W��e�R y�k ���#w��@R�����=0�@O^c	���q�_h_XV]�j`@�P��S�W� �F��B�u��LP�2<�s��Եۆ�r�Z��?B����xf����(�;\Q�H�"�J�*��l��k�v,~��]h��p"xy)���1����)~���׼��ծp�)e�!P�Z�e��vbjZQ�=U m �U}z����}W�Z5���՟���n���PM����������}f�m6Iy�&���r���H��A�&��Ҽ�����/�Ο']�@i+����a���%���ҵ�67�#ӑ �a����-�ϼ�E�[0+$ok[�����SZFf�vޮ����N����|��;Z�LJޙM9A�$\Te����'��]cQ��.�w��';H%�&}��mp#��"6- �	{ZY]SC�r��9��)�}��ɿN���W�B�<쇖i�sn��ųN�3H��Qo��w���œL�m��IW|`߫O����4p��z'xn��k!����LzzC��� �L��~�g�kX��џ�)$��~g�L����ͦt��p[6`������p(�����p�LZ�GO��c؏���	��&Y�S����bH�|݌GR��� �2��l�=��0Q����s��s2����!r]�.�����/u�la	��~Qwy���C/ur����Jf�"X����T�\ns����)���qˡ|�k���Gc����A "�{˨�ܯ�q�&�7Z�	B�;4���'�ޗ�o�����s�ly��­k��XPg\���C��)�� ҫi����p��vQc�\G����&]�Y�_V���L���I*(PJi&�$���X���osS���?	"~?�Xl�ݔʘ�E*���Ɨ�%}�Pt�
���;�{�����x�)S�f�Z��՟���D)����������G��do^��MZ�U��}1(gUB�A4�+��@""��ʆ_P�r�^�0B�ΠY��t�!k���	DD�<} �:�����.��FGl�?�*�����;y~�G�h�AX���1���.���ړ�HBLL1C�;��<,~e��ɻ�[T�#`C���tV�Ⲳ�>��Bo7�P�vc������ @��z����zG���N�vD���Ì�w).���}ʈ����n�l�{�ڻ�4x�I��>�п��2����Q~մoʳ<u�̓{/L��1�»���c��/��� ��E��ڙb��U������3��WgW�w�c��,VE�\F�ځ�� t�-j�#3v��<Oc�*�//����+$ld��%U��9���أ���^4��󘨞�zR%���)Z{s�g� ��=ɞ��j6�ݔ}Q�y
VM^��zW��l˪TgP������e�D��p �?��;���ο/r��S���˷�c��^#��O����߾�qo���Rq�H��}飄��4���ի��_���"�z~Y�;+��<���XSvW1q���11߷��dh^^�?}P=��N�����'^PD��h`����֯��߹�����.~U<s���b.�gE�!�e��XB��)̨:���>T��
��m߂.g�E�~1�}_9��7�.,Q33��0olA��%u�=/�C�}_��Q;
K�TTW����Auk<:&xZ��/gY/Pec-F@65�|$G���M"x�Q!����99�NMi�s�n�K�醱����<bٜm�E�z��3��B�b�ȓ�Q	��B���*C{ �$/�̼�S�R��e�l�f��P��ܲ�:�/���eWƀȓ��������A�0S߳<�2C������8fi�,`���"""e���c �.����2� �&>�~U�������a�	����A ]Mss�j���m(�$����T��$<:pPm�#N��}z��f����PJIu��� ���7�~k��`��Za	٤]h�XF1��L9Y�˭���R�R�?�$M�~�Ӱ7����+y�z,��?�O}qm�CsHZ �~�O��B�����n�Op�o����m�SP�_�0q%=W265�|�\&��J�����e������,I �B�k���)��.�:�ƌ�-����b�����hFPM慨����6�d���o���b|a��mK��Ni��M�{�<��gw���a�[��_W4I��q��,�{b|�#��5���
�q3$��9{��Vl����m�������鎟��MA@rs�Q��"R]�l�Qw��~�:���xIz����VǬ�j�Z|�i�
kYe��` i����Z5�M�B�(�iy�V�њR:�]�櫲����p��UF|�g�6(��5�l��3iG�A�!CI�y�1�At�2wukJ�A����}����)��<Ǘ�����r�/����Hz�e8��B��?�1>j���}I���7%������X8���bT>���qom8�q~A�Kt�c�����nnn�Ye�W���MV^OY��i/p�e#Ǔe$�_h���K�Y�3�9���tgZuoߍ�����L!Y��3����mrrp����	�6�a�J:��������ML��b�>_V�k��Ɗ{�EN�J�F��Y	��`-�/>շc0~nL����	U�ki��Iǿ�n�i�'�E�sO`��+~0۲j�~�M����^�b���ӂ��L��`�]'�F��A��$q�'���\�0����e]}�3����+�D�Ԓ,߇�\���B��m**+�0�Z�ڮk>BATc&X<SS����C�Ы�ҏ�~*��}����ɗ݃�6y��������W|%ӊ�u�!B�N|�<3�g�����y�Vn��{O�Y��̞�(�g�L�P~
��6���������M$���*�3/A��5�W`�}3>�����,/[d�*��s�Cr766v��>lk���L(�'"J�l<�}A�Ь�� ���7`b8����m��x@�dwFÛ7���	(�o@��b�[;��,����"$�2AOo��]��D��ֽ�������r���kI;X�`�r��L*a�)�G�u���GĴy��I�c3�Y�Ĵ�쟍���F��} T��)��O���r;�.��/�=�5��|(zނu����	��%~����k10�n,Cus*lh�AC������~d����^6.�?���.'��hzz�p|�=���0��`��6�br^�*��@`�E`��y�ዯ���)^�뱑_�-H�@�˫ˣ�ƹ"�uuO��ύx�<��+x�M�kg0Ǐ礤D�ၣH��c1988FFG#Rٸ����`��6��hM�;;^�ď~0�!H�	P����1v��,��T4�3��g��kO��;���448{����dL�,�������,��A-C�T�O�Lr/���k�2����+Zh[��lxylȱ�xc�*��{y��@�iލK@�gMOVƹ83ѣv�c�\g3�3ǒy�jdeBTدr���*���E<����n
�@^-�fc�����q�х>�T�Ԕ�ǌ�{]��(99e���My+**Q����~@�6�Q<��Z���TՋ�4T���Tt�eRo�3�r�����G���8|����y���$��
v���V�B�C)㐔�@0,�y�O5�d�Ƈ��c 
$!r�W<�R;��l��u�ͭۧ�/|�y��)����;(�*�mB/��(䯗�߼r��X6�&��V���io,}���	M��ǗF�^����8��QE4�7>��GY�D�,֨�ʁ����_��B*M�J�� 4���q��(�V�M;c��e�SIiJV���e�1 !j���-��������B�t�uT��jN���]7����A���$*@�Ę���\˸��+R��b��HH��3�sӂ���5����^|�TT�nhV�T�ђ���V�i��<?X���#��X�R('�_LC�
��Q����T��.�'��9SsC�p�����=�ኺ�q���-:Q��>j�!z���(�=�E��F�ѣw1�!���~�����֬,��r�>�<�>��;Ǌ�v�Vc����E�w��7�_B6��76��&�mn�t����r/ǅ���!�:~�p\h����E���`�%*N�p3}��ߟ�)	ro�]&�rrr� �20��F���z��Jz*�Ta�J�]_g����LƮ��~����ȧ���o<�/��E�\�i��dl��󓏻u�{�uT4��rM-ON�Q�Ut[�5�0���t~0}X�An��Wg�~I�*d�h1,�u����[�T���2>b��┬&K��vksX�TO@�7�R�k��M��UK�`{2}���@���P��U��@wZ5�E����d�Xq/�;}�z�zY�Rn�E���1�?sV�UTT�����d��e�¸���c߿[o��M6`��g:25H���G�I�:���aj+X���x�w�BP^��,P*��&sPKSZZ�}==�'W�XW>G�0�q����V~g��/�>�f�C���Rgg\\�xevmz��Hּ�Y�e�d�z(������&�+�y����Y%�Y��dԍz�SA���l}�l�]����&(H��<x�~x����U�=������������CKK�<�)����nhP��=�+�H��٢2o�-��f�0�ۀq���b:��^�h�DIb���K
�E~����Zh*�f,�-�Z>\(gz�!�B� L���'��n��>�$��.v��IJ�p�s2p��#���Ӕ*��/�`��,�w=JE:<O{>+�
���Bb���HqCS��4�^D�ϛx�zY�����LY�Ř�B���<###�4/Lĺ�R����/ʷ���h!h�v��:#����9�*-,�S�����s�ȿ���!{�j�ۦԷ(� I&�+�{Ǳ��per���p��#�49�"�
ۣ�KNp=�Լ����u��Wq��{i�{�4����۳<[����������49ID1oݺ�������~i{��� ć�nR]�]�*�����R��%ug�f:�1��ݮ;�O���o+vw�j Xh�K&�:�����#��w!���0�D�H��k�tXU�ɤ����^�3��5-;�ͭ�݊�O!��ta���]���s�5����f��K�y�o�6Y��˸.c��}I�vv,5�P��?�_�$�cD���Ц�9��Q"1ݷZ��@q:��2"mΒ�w:_�g��hy�&���=��D�<��<�7�����d"�߉�
�_��Z�/l�y(-�j�u3��܎��P:��t$�6��Rsf=C��0݇�x�@�������:���J�M��y)90Z�0[�TlO<���U,��% /-C�t.���¨&�oa���wq����Ķ`Z�p��=��6�kQ���E���ѱ� +���`�!gedpt���Iw�07�+�;�83#}���w����qZ����p���ޮ�I�:�}�H娎���l�]2������qS�����1Z#S"*3�	,����e�:ʟ���rKR^l��� S�;N>�J8���!������m�����Ƥ�!��E��׀է���9sC�����TH�k!��^e�G�E�˞r^-Pd �ڦ�?��Bv8�ʛ�c��+Ыj�|�G@�3��JQwjb��㲪�"���=�������~>>B�d=[[[2��ƒ�I���+��!������#��&3A�1�Z����<���P�?�C3��f��R�Uu��߲�L��Er1�"	0KHq]PB��W�tA��4��$=m�:^�Z���7;�I��ԣ��
-�F��w����:]�H�ۤr�=f.�J�'[?t��ʔ�0Q�_�{dP��+~���EV��y�oVw�e�h���|Bd����(3��[��g���X�ٳ�z��^1��Y|�{7A	���G�O~��ܫW� R���T���<oT�t�r}���T�3?��\YV��Ҹ�[��V�M�0��� q�7_G!���^5�C��ɩ<�i�M�AK=�m�]0%־.������NM��Y�`��(�8:�����m!C�˿[MM�V����pE��?�3 ��`KY�V���y Tޓ�XF��*WN�`6*N�XMx5�;�Î�z߷c�d�jeʽ&�?H���f
7�|R����|Thߋ�{��I��
���?E����qldD��M�"�_�}J�?�=�*.�Cߍ�����/^��Ոs�[��~���.��o��e���Yp�7В{aW�U*,�!�8K��C��B���	G�&&A"b\e9OO��8�D\\\��%͉z�q��c����v	��l�I�����6a����v�&�ҎM�?a
�t{�<��������['���<T�db,flllh����bz�ĥ����}q?��Ub��^�I,�ղ���Ź�+�1
s�N�#m���Iiw����
�:N���L�R����V23z榚#0t��� >I�xlG����g��OeTf�����U����Z���wҶ�u��-�^=<<��R���t~ᠵ0y�db�+`fu��ڽ�Y�2q�0�w�ƐFQ���E��vLgh�Y�R�9ʮx�$�9�f �&�:�� 戕��`}X�%���G�jk�&���f&�%�������T������@E$������&�B���^x�}X}�6L���=�T�m_U�8����Ӵ��Jm���M�Y��� f��k���hv��%�y��m7n�ӶI��쉋����Ÿ,���dP��������@{e���P����'-dN���ę_ 0�+�y)	V�:�	yę�S��6�잏����i?�ܚ�\/,nE%VT�[yZ���~�����p&�$�\�0E/���k��g�7�m�V��?�3����-��*�w�m�O v��w�z��<5{�P��T���SՋ���r�K���n�/V��_4�Q�N�lmMm�H�\Z0�t�L-��hG�>�r��}ʕ�J���h�b-5-S��XrJ:C�`��j�Y�Lc�f�����"����0~�zź�稹ȝ3�$���L���M�����W*~��g�����_fD��$���l $  ����� �|������m1&u3!<;g���Hk�����^���N�{���YV��.��E�n�X����
S�b�*_�k�������������X%��G���_��,Br�d�7�-���m�t�7�T���@T�����z���Γu�#�E��&����=s=��ɽ/"��!�`UM#=WϜp��ݼz ���E�f Q�	 ɘ�?����uY>����sW��^aa�hs3�>ߋ���� �[�;9����D!K0N��.d.��4|,Q'TNkˇ�L��T���'��1'���B������C�p8h�n�G��^=?z��]�Lڰfm.+#
��<v}B���B������t{Sp7���t'u)��%2%��p�u��cPʃc%'�����6� ��Y!z���'��2��ܺ�ɶQa�����^CH�*޽��勖�Q�m�q�a&>z�H���Ȓ�8���_h�6�SM9���/��ɐ��������!����p-�����5ϵ��֐��@v�Z��^�w*�����k��3�=���c�VVV���x��LP�׋\���J��P�o�}Ű�3��fg~��I����f*!q�*�/}����(�W�-�)����˗�=�E�Q}�ݼ�h6��؀�8h����!�6I��l��mW�����`���2�4?��!b���������@g�N:��,����Θ$�����jUkkB����%#�/��KAL:>�+�&S�D��t_YnW芐�<� �8p��X16�H�O`���HϠ):4ee�u{E�)ԍ�U6�����r]���Af���+yi/bn�����|�KGGg�Ri�$L���×P�l��g
 f��c@�>�q	LˌIk@�̎,���%Ҹ��d>wR��\���	�_��Z��0Z\���귉?�+�2��Q����yd(�&/�����d(Հ�,���}C�7_�WT��.--����E����w�U_잤̬��H>;�~v>etR@�B�����Z=n�޿�-o6�����+1�:#֔�#3��?��%i,g�c�TS,��߼���h5������;���Q�\���$��V�SX��%F�k	t��I~�K���|~xmh������Ygv�๟J::~f�e� �q�;�Ι(�᭛G����%iH��n����V9��`��y���v��j�s�:�}T�4DĿv�������]���W�&q�qu����<��-�r�y]��VVl"N����$����4�M���`��I&?Z��];Ht��f\��dQAJ�E�Bb�Q9��K�����;?�����6ﺻ�,w�$%�ë���"��Ƕz�Ȁ!)�;��Xi�9���� �m�g+L�Z �P��՚p������˧p��F��z�{��+i6�+`N푷�2�][���eg�f,���G��0i�{�y����b흓Bgo�P��/�F�|�%D�j�WH#�D5�s+Z� ��b���zǙ��������1���m�:�F���|/S)/-%$A1ZǄI�
F�.�Rf?.������,.� ���&��N-�y�Ue��Z(���x���=��FmN郎���n���}�ϸu�E�!K�Jn1���|����H��q���c��N���؀`����:3�d�[���
z����������	ε�i�
ђD�^_9��s��Y�3�V��[�~�9�I�Ϟ���+i'VN�H�[��&�)�_`�џ�]��l%��v�x2�1��{�/�8f�1;�u�f6���j��=ײ���_5?f�4l����UU�@!b-���Y�^+��4�=]d����~��iP�Asj�}-P��G	�C�P�x��~fy�����(>e�����'����u�ق��K�^曒�^b��ܩ��K?���t�m`a��I���c�K!��h���XVq�:����}�vNX���%f�c�	�F#��A��M��cNX�D#J,n��B���h��G �9]�� .S�KH-���o{���]qU��D�b����E_�1���y�v���L`�NA�dZ�o=�7(�}ΐ:怳�|̼�P��b<����� k��
H��:o�#}�ɼT��٥
����>�Yˍ>%��$u�����Z/Yu���|=Q�a����Fl��W���kAF�f��,��X�Y$!Q(B$LY�dp��e�>D�~��i !".��h.���A��c\�f�00�`��~�|̿9��l���.�+��vv������h��(�����Ȯ*��E������y���U�<Ą�3՝�Y!��IQv���C�����_�~�~�'ר��>��E�D�P Ʀ*^������)��"���ӈo
���1�+�(	-��]�;��>h>�RMm�wsN�Q6WiP` �M���\&�`mԄ���ߋ1#����Q����kD���<���I��lV����f,�d���G�z���֥G�1�K)�]o)�j� KF���7W
���S����^\�����$VN�-l���.�!�����	p3��H۠P5;/�)���GC8H/�������;%6^^�oI<b^��o�["��k��Ѭ�9�ˤ��1�,���U����jl��h/*G����ѥ�?jQ9	#Q��n�'ăS��%����9���kw�h���c��B�r�K��w��Bb�0�ۖb...xX��o�o��h�P������S+4_m���S����YI�~�0�0~���o�?	
��62#<x�g���Bʐ��`�@m޺V�s�m������ ��2~Y��#�Ct�],]{��R��힦�4~�󾭬�h(@��d���.�$
@@���%F0���Ő��0�ŋ�D��b�gk�߼��:�e��xJ?0��}}��<���嫪�5֝y4�@~�4p��;".�*�<-tl�����Y�+���E�'����R�u���Q~���*����������T�X�h�E5���]ʪQ�? �kȸ�4��p�s@7�������˘\a[��'fz��LN�(Α�F��J�)K!X0��1k	ׇ'����{�?N�vۄ�Ӗ� �Gx�%��J���#�tZVg�����sýi�PyD�r��V,���k#xT�A���Xg+�����$	�om��VA�K'GJ$�4�hm$Ga߻9�@d���o��*�;7Bʊ���Bl�_��8�X%���X􋳲aG���vM+�p�����ϭ���=&����5��{I�z�O�)������Ʌ�?��+��d�n�mll,"�ڞÚ_X���'{�tYh��19�(�������>4Z�ؘ>w��j�f"�����گj��(�r�u�a6LUA�n{�Zz���z�Ů��y�y�����aL� ���� �B�1��o{J�{R��@��ppr~������E��Y]�r�<wg��E��T�*�a�{{{�镭�A&_ˡ��u���뭜�I�2M"��]�|o)�Q��?�}���P����v�V2u��y	�`���a
OAs���9�h,�S��Z���l�"*��ل��q�}��-)
��<�ϭ׮�cڂ�7l���E��4B�L�y�?��9���z���_M���t��d�Xো8�m;�5E��`��wve�����*��7W�Z�	�v��d�� B�x��$$�htT�q�+�z��6(�e!k���N�L7'aׯ����i�dl=��ܕe�Wn\��Q3bWb�� ?.�A��T!���Y��򊂫���`y���Ґ�|�H�4?�,�{�#����7�CcWL��G�Z<O�~����V]/c�et�#��ӧ�	�����r�\�"��K.�O-�'b��]�iG~�51Eu�;�:llh����M��=	���5����ֿ�#��0��_���v�U2�e=�h)s����vjR�����d�F��=	�4Q�Ԁ,�fݓ7�ݹ޾�� d���EW�w�k��}Q%��o���w��Hs�L�Mv7'�m�!O�����k�0�۰�aL�����R0���Φ�?�mԃ|�υ���GV�Z��F-{�9��+����:
̿��ׯ����u�`����)��%��Ĳ�5�0bo��m},����W28}���c
+�0�T�&ezd�G�t*�jŕ��K/�m/!��iYH�p���*�F�O����B�Y���W������s`x���:b����G�K\p8|�Ag���N�䔨�Pha��3$����H%$'GQ�_>�^�}��ݯ��BC�����l}�1��v� �8�7!�x�a�l��p�����{8II��%�^�U[��>p��.��1��O'9�\?0ܫ����і�"���+,"��xG��[� �6ƹbn�۔�=�g+.�q��L����	��J36�j���~�TYY���u��Ź��;��� �0yl�Fr�J#Ŏ��<1�U1�j��GVc��q�"Wt��6����ӑ�]���s�:jHi�a:r��Rtcrp�W���-��|��=�K�9�/_��6����)���`���o]z���V����N�/�{�y>Y��Ŗ#S�{��C�9��������u��d���P|���x�7��`�(��)��r�R^jj*Y���-��5��ʧ�a3�xL�C�V���Q�O�����价����aQd�/�d�7�ۧ�5�J	7.8����Tc�>cD���<*{o� �\5�}��F�s��- O�o_@2�,�P9�пKS��;G����c�a��¥�6�)���2�?���*�F�N;��3�>ƅ
��k�'�{�'=�����l8K�+��)��S����C�m"P��ۈ�Xb�*����8�.���;��kn��nKl?ũ�t��ws��#��M��4�/��faq�jNq����ʄ����Z]�N�4'0{� ��L�L/N�����Ɩi�r�f~�<�>��}����8|e���VK뚰 �k���$��Z#...X���'=}������f��9<
�9+� +�)$���t�%=){�3S_ҳ ���I��֕k��c�[=%U��/֯�#�w>�5\�ՆD��&��_�9����])��/�mC���<�K^��]I+�o?�x!|��Wb1bq�9�M�W!8t-�Ǫ��AII�:l./��}�)���y��+���qG�u�aG�%t�������u� �z�
yǮIZ�>�>�3��3�h���{��5�2��|����<|^[������w;�E����w����v�؃|�'��d�n1�=ӀB���y��	�|����}�#	P����`Y�~w��suuQ.j�\&�T����7;O��B�C�*���:�zϫJ��F8~�<JGȭ|�W�R�J��`�ܞ�0ͨJ��,��[wZ=^�Q�Z��?��E�4�P;�bw%�T���I�P�f��q��eAH������jf��T8����m����E��%���ˆ��A��7_�,z+u��}�5ꆳ��5?D>��#q���;??�N���\��Pȋ�n��A��D}!E�`c�����D����̘�`�� �*Z�L�F%2��&ӽ~���f6�E=�֜��2��F��g&�5a���}�r������U)��!1��y�S�By�^X3f��m{�n�po��S�8"!O��M���]����~����P3����l����;�������+h�7.=3d#��=��A���kjX�0��X��}�����~��_-������b�-�.y�KfR�6ˇ� III��H\�UN"s�RD��`z������fn+B�\\��#�m�y�p��Ǥ6C�q�bP~>�\������i�JV�E)����ؙ�ؘǏW���-N�cj�-���g�J�f���Y�I;i=2����9'�Zk�gxX߻ƪ�ݝ��q.t�e���n������;�[h�u1xJv�ǯ; �y�.��D���[9������S#�,&���龖���9��PL)Ӌ�s�oݺ�f:r�Ѐ�V�>X�`�a ��5Ǒ:�vж�a�����~,�||u(����V�4�� ?y���6=�!��*F�
���j��b_Au��K@�1III��(2d΋&�!r��  v���|,�!$�P]��P�}���ygQ�,4�������|~R��f��U��h*ca������;{H�����; p�e����vG��9���n~�(^w������ֱvm0QVW�/�.�+���׀�stNF�:u����'����r����M"I厇���!��$K��C�r����H�<�_�Oo����»~t��gg�>7Ou.M���j|C��_��L��w�a���E�/*XE�|�_rom�&����6fy�n~�R})9JMn+�>`�~z�o���ۈ��� ��Qz���� ;��lSy��������6��d��̨.��%k�B9����m~z���Sy���UG ��L�k`B����� 0��ě���]�*�'I�7=�O��	V��)ij}��U�s()M��ø)nP������y�_'���Z��[�H�z#�ݨ��q��5*}Wa��m�2�T u4��g~����_P�SZ#�����ͭ�fge~ ������'�%����uܗĢ�eR��"7�ǟx�_�#},��=�*;a]	�2}c���MW���<< �yX�l�9�NU::t�A�鿖g����;?J��;��a)���MG���U"/ȉ��η4���A����i�U
T~��?�� :��
,��[��ld����F�@__?��,L�q}����[�jL-W��Ƽ�X�gn2�mc���q��{���/��45{�q3���za�=C�"N�8V֜�(T��V����Q;n׿��[-�	E�>�YTY�r|C���w��E��iꚼS���p^��5�v[�[��h5��GW-�i�_=��� II���;�M�҉	�'�����͍G��g����$=蓯XϏ/����������>. �E߀>UY���|�� ���VдωAg�&��T�~��G���#nL�|��zA�/������P(�DF�M�)��nn�sZ��Г7�@OO'?f��Bvs�a!��'IO|Bl�*!��['˂�:<|�0
�d�n��ģ��UKnJ��oo�����O����k)�4TU�T�	Dd�
6�.�3��f�X�^�}�2��k�����57?����5����z~�g7!���+۬ ���_�ۆ�>�� �J�5�j'HRb������v���`���Ƅ���eM�gG��FÁg+����5c	+pSz�/H�\��5�y�5F�,q����v���{r�������4�OF>o��c>x�X��]0�I}�
b���������(W�9]���0�s�����|OR�)��:�jQG�a�y��36�D(�6����8�@F�(z�1£�׋ftm@�:s�#�:{��9�V+ȅ���|��G��E��%!đ�>��Md����Rs����l&fi�^�O�[�,�ށ��V�̌���@S�(|�ޅ"mP|�X�a0���������2������NwǪ��ךd�zX�����r�����z���2+G5_��y���jx���<+�������T<��:y��Kc#*!9��s�v���v�@T?,Uͺ�xU��fnaa��'����BI 6"��~�����ҒYb��� DPY�����6�.�v���pR#���4�}}�sBv5�������.:��)oݰ�Q��)�O�0J����o�M��ؔ����.X�{�Pyj���~(i1o��N�4/���(�d)[c��(|�ʑ�xҾV��͹�s�*�s	��+�dB��)2*�bl`C]+�u�x!�<�Vsv3<:��<�ĄLk׀r��0����0&?$6l�今������ʘ⻸��~�*l1��])���ǵ^�T��`x�`��� �[nCӥ�:��\������mc���uqt��c�a�ͱ]���/����~��5R���$�r�������Ԑ>`?Y������_e�
��T��Zp"޺#��"����W{��>f��Ԃ���rP(U0��^u��GS��T�C�nʂ����]�-(p�ۭ�qm��ycv������-2���_�k��}� ��ڍf���Vw�s�������I���Y�2�W�l����Q��Y~�w�,/���)
x࿓;���rr��ŊOJR���u?Z�44�FQ��q�,!#H�ivsF��טx)�Y�<Ɏ�֔4E��z�1\ R�g��3p�G�yEȷ�8�h�R:�M���$��^�h�b������D�b?��cE:����V��-]m�)(��X����?ʍGG���hc��e�o`���4�7�܏�����U�r��P�lU�ʁ]\�/N���l�Z���Nw}y�������ҁnv����������99�k�����j:�=���f�������>N�\�?r�~ {PR�L��0�p,Y�-V�ě��b]�Z[r�23�=��C={�}j,'q\�MS:���?��7�9��z_�������J��eT��W�Z�[8L�F����xe������|��� `��
.WT�Z6��,`�ٹ9Mm�h���$�~���9U����d���d�;`�&�:��BK�Y%O&�;��D�5~:`7+gS\�_݈7w�����i���T�WL�k:�
�I]�+�4���=�Z�k[G�t��U�������xo����w.�<�#�,��@��YƩ3�X�>uuuʪj�Y�ؗr��+T���O�������=�uT��لx�e�����X�����Q������\���=<=�Hm�)�rw)�[jv��F�&�t�{&޺�|�h��_~s��
"�ҩy���J���u����ǣ$��������04 ��S�w�#�d�j��+��*������kg���O>y��HCT�����H=�zW�~�ͺ`�բ?���A�6�4ֆ�+Wkܘ�rݼOx4�v����7z7!�e�R.�ԯ��3J}��p�K�����R���?������Ga��֜�iab����`ئoh(���.�_�xT
��E��1��0�����D����N����e`��2}��#X�DX�f��P?��|��	)%e�(�.�s�rs���)11��HƄ ��F�q\�E5v��Ub�*��ߣU����ҡ�ѵV�,/W��L>,�6�w��0P�HP�J��K��k$d$C(H7������iyC��oM��ٗ��m^�ê��������|y����8y���B��{}=_vGQ���鯥��8m�O)��T'v�8�]�*v�O}�4a���>cV�4=�=�m���� C>̏k0�u�uO��ӷ��**H�G9�������"����DW���o�^�7���{�;��0������L����܆���"���nf��6Ew$`��$,��f1�{������AG|�X�:q��-���B��,��#6qڙ&ϟ|�˗^KZ���d�	�>�q��u�U�F�P��uv��Mqp�w�`b�ދ���*(�~�dYX;a���X�y����� ��
���ut �WT��#e誷	˄�k�Y��E,� h���uk�)���i�G!�Q0�z�έ�m�ȃT_�b0.����3�ЇB������n����4�̞�����[8~�S�Nv���υ�w*�$�N��?t�ȟ�3�w���n8;��YLm��S����`��\[�%�G�8�x�a a�PcL/���^���u-}�ʛ��먞=�%���y�gyʵ�3�윕X�dܣjz&h�-��Ekۃ��8�M�X�5Q�Qz䞤�:����--��'x����b�)�������9���f���F��BdY�,\�ml^V���Y����o�S+4�o�m�X^�����H=c�αX�Yh��u�WW���v��W���ٽ}��ߟ�q�-8�~t2.K| n�>��l
�)6=�E�}x��۞�bmm��gpkR���B4D4Lt��6���&��p�j�Q{��D ,�f���MMϠ09��u�--)[�p�5�@���O4` ���0j�03�i{��Q.��ܐX���������3g�g���
o���o��,9� �4�����4��Ԥ�~Y��Z|�㾯7?�"��Zs�?�՟��tء�
���O�����/c�|c��p*0F��- ���g�o�&5&���|�</77�Y��R�~�}��T�Al!��R�΍� ���v'� )u����F=�N���L�Nm3u�ԏ!Gg�f�S�*}����wn<^�U�6n� y��x��F����B}��p����LV��m�����h�vڒ	7���z�x���:R���+���V����iMM�k#�۸?�gD�_���'O¢��_���i��SSÖ��\ZJ���Q����z��s�'���N�I��k�ט{�[/�?�\��b�����ͺ�8�ڞ;�B�T��hߟ���\�h�Q<��>3?�I�cbUTV޼���������3<U����?�v~o���
z��J||dD$$B��`�	� ���H���$�  ��c�������y���D��3��Z��Q��������~~Dv�t^4�XY	�Ӝ]hh`$f����;$�1���sw:X�ΰ�c/�h�hx���N���d�D�m�ly��(��&���j�-�Lo{����4�R�^�_6�*\��cN�-����m!�~'����,*m/�e�s�R �� Wo�����r�r�%��ݛ�
	��;�Zնݨ��|#!,��*�ន�O����K���D���2 st�ɓd>�ʇ�����zw]�w<;S������;р��%^���]�--/4=q��f���W���ܫ����y��i�f���Pi��=eu0Ɓ����f������x1���� �u�В�N��ҷ���a�����K=���V�G4u��.�oX��J��p�P'r��xV��Q�E�y�Q��]��v< @(�!��>
P�5���z��c
\uk:�R�e*~��Z�o@/�&''�k�t ���m��`��O��3c�G�ڂR�{�� ��bՆ�F������޾�4ΠҬ}���s�x�X���Q
�]W����DW!�����l�R��k�c�ڪ���2}]�$xI\vE��
"���܆��}dJr��.j��8֡�H��*�-���5U�'� �Mbbb��rɄ�K]}����Bz��T�c^:��̈́'��y-�����3V�ir�NP�4Mt���(111I/)&�{���Jy���m���ȹgN��|�s.��x�q�Qy�q��/]Y6bJ ���ٌ.�f\`�z�!R���*�wĘ�+IW�<��3v0�9��T�jW�U��#�aG�p[�v�kh��6��+�q�|�{�f��X�d�|Lo�%
��%sv�#R����� �j�a�FZf�v�[��go޼�אP+������V�>�&lj�c�lE	���5n@3pt�j�k>����ɖx�v1��w��������2/�	���E ²��ɋt!(�_x5��lzp?���Ʋs������SjHl����#��?�se@^z��̼�f"���[��s�]ĞM}̮�>｛���X�P��4 ��k
���5��͙yyU�,�6��D	c�=nӕ{@�����W{����i�H�@�v:r��/�Y��J���^���U K�lx��e�~!N5(��t%��Y���Ńݼu �R��&�p|���������Ε���2��"	V��^j����&��^�2T.��x	�:��Xy ��E�d#�w`�5��_�9�M�ƺ8����F)#Ɔ^sڳ"}���?����7����E��OX$D����<u�x����WY��N#2��v#��V���m�&��� m�ܥ��A�d�ߎ����F���n燧�vv�ԈlD��,i`ᯈ�ϸ�>��`�뺳��	J��#�u�2n� ��E�_�ǼUX;hc�gM���	��'�������?~�OcY�U���.����>�� �a�Rգ|��	���\b�S�+�N�T0-,,�R�.60����C�,�d/_��W�q���+�4c�#['�<0c��,3�L�[��9`i��^ˇ��suq^K����L���Vt�u*�����Kn�3�&(O☔9�Ӎ�gtDx��faVvKK�n��>��6���b]U��yۏ&.��tf��A��A"��JحU�9��0�e�����±	�|�=�L����/lD|���Az��@�k�U����?�CNa�c�5◐X��V.����ʛ��M��.���㭃�z�ƪ�t���K�q)�]�1��cΤ���q)L��_���L�v��L0�� �cO�����E� 6ݦh�}�	+�sas7��U���<o�x�f�S,MM��~&^�ǘ�B�>�{�WUD���c���to�̒B�;|qn<4��Y�-�ȟ��l�a�pV(������X�cln����|��������C� C��9?�?�]�(%H��=�%�{$�š�%��ΐ����0f�/j��W����C�`��]q���ZTt����'�o�6�|�3U���{��F,*�5��V\��D����N�2������u�������݄���� �M�up��B�D�LV���ϐ�����YU�y��Ltuxe���\Oo��9 �oZ~)�׿8��=�C絴��%��Bb�E��	niPTBRF�깎R5ׂ��2(u˸ n7�S]���� UJXͳ�f��5tvNN�f���nns��n�����Vm*G?��s���`���Ro��ƒ�����'c���0�ީsy�̴�cB{F>55��z�W���N�e�S����˗���I<��9�i̽�~�x)��o�����gbrR1���J̓a��CB��ѷt�'Ƚ�bZ���866d
�l�8�����۶/j��P�5�����.{mkq��)f��ԋAҵ��BM����s�������:
��C���ݴ+�\����	9~�Z�}���1f�c�@��Ϲ������@^�qn�Ǘ��5��߿�z�1�F#!�tP���ĥej
,=�CCT�P��)*��{ϒ����Zjjjj�)f��
qLZ�����@���=o�~)�X���=so5E����i���ˏx�����+�jh�~uZ  �\��٥f+���TA6���=`���W�\��S��9�i���!6wG&U8>�eGW?�x2�O�B�{��z�׸J��J��|a��s� �De��ԑ�Q1 W�\P�'�w4�/����+�`w�K�R�)���+ja��=0
B]^��0#��p��,������O]�H.���}�R�s`�Y�uJ'��D��Դچ�;  ����q����r��
=�!���#�N*3��D��a�ë�sֹ�
�<d.~����}��$3k^�����oD�����	��O�v�G��M`���ŵ����~��'��_[z�� �ət1D�\i�,�IF����f&&�z�|����T!,ͻ�BBA��"�+���Rޑ:m�����H����ڶ�`�1�|��i�0`�.�������?�] x׺�4W��Bы\��P�c�**���A��{AZ�����5��7I�n��?��؂��Nw����W��������0�5����n� *�)އFw����SA�f�ܰA��]
����A_�Z��Ӌ���<ൺ��q�S�v���~��ǹ�R��ib=�>����|!�����/�0My5�=Q�$�:U�?�64Ђ�U�5���_ZgKK��W�$�"I��ˎa��j�n��en��7�F8�C-Ķ�ϊ9�G�xU�����}P�
��oIP��9�p��bK'��""%]��}�$	��_0LN. �·��.t^�~\6��VX0�C|	�~��/�;��D��������V�;O��qN?�y��.��$����?<D����T}uXT_�.��"-5t(%�
HI7�"H��0���H*0tJJ�}��{�w���<�xb���^�}�^��	�UP�l��*E�������I}�JTI�T�C�n��[��EDx)^`F�m���î�!c��k��T� �ü��pa��|}%��_�LLҤ�~�8
a����{�����GF��si`J��( ժʸ:��G@�K {&����r���F@rZ+ɼ�T \�cx0ڰw�wd�,=a����%Ԙ���10ss{����jij*yx�V���� ТC��COL�NG���͂�Ɩ���%��%r4�rWD�h�����6uoxz.����*�ڇ�q%�w�����x�=agv��_�����t���r"n�nPз��Qe�D�g��8O!`���#W a�onʻ	�W��~�a��";rde=VP���W6j�7�S�k�ޡ�!���i�okƢ�́��u~Pa� ��.2qwl�Q��@U��;ז*��r�wB�Բm�#&i���~����(�iМ�Hl��u�۹Z�I��Y�=ϻ���.4���f/p�UV�{����x�]��l7��0�+\��M�kWP��w+9���=��6y/����4؁k�+� �_���i8��{�8%�ԫ�=>�>W��ʊ֠)L�B%� �aaař���������~�i���n�{����O�u�eQ����y�a�Ρwn���?���}�飂��T�Yc �Ч���C	�Y1�m���s���]�@N[{r>>��X�,$�x&�%m���iii����a���3x����.�����{_�k��_�&*E)2�ގ�T[.wc�{�G�i���j���\^�7:ϡ!2���U[�oo����;�����Ƹ�5�������ӟw�n�Ǽ�/O�uU휳@����o����8�}d��7gr�-&��br[}Hm�y�m��S�ң���n���4:_Ѷz$<�gó��%bؖ�X���-(��%��B �݌��I�6�5XȻ�2������e���'q�!��>�B=����#��+Hff�'˦	�С�g F�B���1�)USy�
�LKS��6DvK+,*�C�Ӛ��������S�t ƀ��x�*�7:
zb�qs>({+�'I�Q݊�\׽��k�_@*�Vz���3���S{eeB�I�i_���{�4�`�*'����^=XQ���9���}F$�<�A(�O�Z���Q�G!�]���I������Г����g�P����ڣ�_�m���}�7^~�k7$����q��;ʸ��E:�΢�S�F�sCv�W7�[������ّ�_�̗�9�[9񯳺BWQ���I'*y�AD�F69��Brzq�������k�)o/��k&gІDl���5
�d� ښ�����wN�7X���zB~��'Ѕ������:�,�b�Rf�A2�������YX��hr�s�5 �wGG��������z�>쪵��HO�� zb����o������[kFl?�Y�d�VGv�Ev��㨤��:N��B%/�ԏ�J���P'>~�VB �*�������
�8X��-�Ehhpp���+��l��!�����^^�X��	�q��k�RQ���G>�F���p���)���eٰ�MrrrOs� �ջ!ʣ�]o�o�xH�&Y�$��Ǝ���O���C3�Mz&\���`�@M-ܾ�A��$�����j۱&����7kAT�L��;tl"҂����T�а�߀4D�����^��0ڋg���u�b{���:��mD����ǘͿ�Z����*��b0׍�nf��Z���`l�P#�J�:���pڙ�Xs�5�Y�ca��8��k��O$�w�[�iΦ���?�2U���l(�¥���M�\��|N�I6�7�t;�sQ�պ����s���!�ɶ,�Vԉ�f�_�e�UNB�)�����o�*���**��+k��ee[P���Y?�34�Xȃr�����H*� �aCҊYX^��c���:VP(���7�aeuEeM��\��Fϰ��)��l� [2 ��p�j�l��x�<?�J��g/k��O��	����nm�+hv�_�K#�J'��5&?k�I#����_q�KXK�R'*;���_�����m��:O�~�4��i%ITB6�q��8-620X�:��E�L���x��n��Ͷ�^��`��e?2��<fY��ۢ�!��5y��ڮ�Ohk:�۴889=nΫ0�nn�r��Xf/_K��꫷'�o?X���:¡�2l��	P�j��F����!���W籦���dX�К���f�%˦^��(��ףi��3V���� ��/� �=�fff�$��g�K�Co�T�j��p+�����x�%�'���-��mR��p8hл�� ww��D`(�~�4ll����%1�;��1���.�O��? �a�~k�bq����'#�����������(��`CQ3K~�a����Mn�l+t(�y6���9�KCi���T��
J��������5���
i�a��Sj`�#Yx�)���p|uj�� �)�W��o߾UQ�U,�`��L�DG��n�fa9⯡QU���r��m|�t�� ���!��J����T�d����̱Y��Sdr�J�p(;�j��ᆥ��VZ-̹�8+7)yyZ����2�O�V�P�l����<B��Vs	�d�Le�Ǥe�����
��E:����r��pi)����;n����-�[vy��/BC;��}�@�R�zP͇�͇��_$P�A���]V�J��:�Q8;Wp?�o<�o �ބ��7����ΫWq��)�d���]2)j|�������f�☊�f�?EdXgA2�t=��sL���EM��
Kpߧ�kŻ
������4�)ᨈ?
e�+"�+'�)���\U�߸�{����6ѷ�E[��w���I�F����؆;��d�Bۥm�G��3 d�=�̓�A��}��"�*=`3}S{_*�BU��8�3ñ����F鼞^�b�ۋ�l�v�f�w�}�0�`�r�������?F�|���.Cz�,���::�QLp����'���4�7�C5AF���)�u�^��y�ÄQ���1^x�^�{�������۹@�++d�Sq�#���jq>^^


j��_�(⇌[��r1:�i|��<�;�Ls�ʩ��ꘙ����M��{�q�0�i@E��ޫi` rs���!�e���<��j�?����Ҽ{�]B|�
/�%x1��r�V�ڜ_<\�����T8:�J����=���C�B/~6�;����y��8@���M�(z-�&x5/��.Ƥ\I����@o��7���?9�rJp"���p�G����"��{���TT�v�~O߯M1�#+ŕ��d(��h�bҮE=���� [�8:9�k���a��a������̌�wq�~��Pu7c��$��
�7��X��#ĲyKT��1�� ��y̞�2�E���*�Y�G�n��K#e�%r�E$F{	B>$�_q3i����GQb$fk���zsl�>����U0@/n<�K�0r�U�O��!�m��*�I�q�۟�
9�7�FA�L ��T�NX��|_x��Y��>�|�d�-#c�8(��,DFh3~B_�Ǐ��7��lқB����޵��_�s>KKf\]՜;�i�?58>��$Zӱ����QDWM(a���A��|	��d�r���d��8!�|��*8X<z���������p4ed^h>�/��})��b�͔�ܙ;w�w8�:�������z�G%�ǵ������w�R"a�4["�
���#�g�������;<����W�)q���'������ @��!�5դP�z����[��ѤJ��Ez�{�/��^��6�w\��Mlw��T��PG��]vǢ!�:������\o�iK#V�"���6m��M������87$w����_���tD������;��w�G��Fq�����qM�շ �m��9JG�?R�
�y�)s�U�H�>�lŠۧ��C$X���u�����칄V���<�NX�2d2����P�� �����n�ҋaYr�9�.�]W�o$=�3�`=�OT:R�t�@�NFdn�
ܹ
8���;����� lC2��C;M��;�é[;���V����r���ߢ�������h��������䱄MB�������ֶ�Ƀ=W�y� \/^�oO�0x�@�Oy���l��Sx�=�����u��r��x���'�R}5�,]-Vd�dW�g��
���~���U�ycd�nO���v�h�W�����4up�p�<��@�������T�O)p�
u����?�9����L{G���	=ϔ�+``c�c<�(̖(�����V`�V�nѓY�OIp.�T(��Y{EUX�g�*Y�肍;��鬰1������с䡎4�P�4S�"���8���%��'��(`��E�.z�ZF;���Vɷ~7�M��Ecc 6�ƎfD��K1��u��|��ɩ>`+ �뛛�5�R�(��+J�d\QQ�D,�*ӟU�%K�~��0D��!�_isno��NV����g76�wjS��4�5��T%��F�z�я���B���xPE���B�~������O��5X���S�\݅,l�(%⌣w�LW��"~7��02�B��1�3�2ν~���w�;�tv���d�;��� �أV1��X+*�[�U�7���[�.��`Xm�8��_�w�	�8"Q�Q����x���8bD#�+Z7��%����22�5s��j�ф�#'uz���~v�c"�f��J�Ϣ�� �dB�ѧМ��í|d ���:��Gx��>�BN�m�ᥠ]^nH=�Hg�~m���?�t��9b+�q�pσ<�'�Y�	�w��fA�g>��a�:��O
�}�ܰZ�Rf�~�#�o��y�U	
|.�Yz墨���ɓ+c�V�q�p ��Gp�@�I�i�}��������6A� T���8CV�R�M������?h���!��CmAf+"�~q���`���F��-`�d��|���mi��c�+hh�O637'�2ī@���q��CL&�⟻��~��V��53'��(5�j$��2����E�k�7ߞp���96���s����Z\���OF�؊T�Ro&$s�iq�S�mT1�������L��Rd^_����%��z|�J�c�az;�O�$�մq8����n���agv����/�t1����J{�S�і� Q��q���J�6͂	P�dU�fr�K��s���W$��8�&����My��'Ox�5�W��nJ���bI���cm�����8X<����˼�_�����$~��xf ��m��Ȣ>1ɓ�c��e@���D~ݪ��XS� ��0ndX�6k����񉊊���)o7#ʦj ��l�n�m|��O�����~3���D����*$M��.�ھ��G����KSNK�����B�2�&�VQ���������d�qz��`hȁs�Z�mK����8=H�%�4++�Z4�S*��LK��P�
@���MZ���E?�tuI=נ>o�y�v9_6�:�0�������e�D�`�@u��x�`����k�j�< X�}�oQ�V|����=p�T�ec眸�#�����Y��G��p@�SQ��BO*��W���..�0Ү��8;h��6!�K���� ��k���0I6����Iuր���''"#$$�=yjb�~ ��|5DYf���^SCkBԻVI�����q���YtSc��m���s����5���Xf�\{�`<fE�Ե+~�����_۫����s?���P���k����ט�"�J�^V�I6�Y�H�F�r��۫(�UFq��='����l^� 5-MI�6s�H��|$ł�������� ��=��Ef��▨]�2w6]\"_�v�!�@����uz����o��<�����6�oX?<�z�'�<��^�����������K�ā����������b�d���=ʳ��~7�'�̛YlZ�7������D�/��NV(w��?>t<���'ͭU���7�R�0c�~�M�>��e,]��͸��.J�����d��g���MN�yn�RcE���,���[h��i~��!$��4�YN5�0���gh�n
�I�}T�k��R5V�BlIT����V_AQ%���^�\������� ���O+	nLL���b4��n]T����%�����7�"[#�>C��-���7�}
� @�,����%�D���8(�P.�Dm��N����?Q�O���U��2�*T� ��EN�/��C�D�r]�V�0�L�A���@�D@K~jZr�����;4�����?;�������fNKk����w{���V#�F�p��ʽ�9�^��}Ҿ\�&�������k�t�ܹ@�s�(��3�C��{�ɦ��3I\K[��TT4U��GQ����`=ߴ)v�q�����/m�L?�;߲w��H]Yn�`�n�����.�#�����J��l��/n��ʫ��;y*��3w�%%�O�G�>�;H���cR8�Ȋa�fD�KtU&$��}���q�sb��'줏ԓ�,���P�"mf_� :����Tg[�
!�7�o�HiEb��B>-�
�qqW6��sG����Ǎ�j���ܔ������+ /�$�x���s��;\$�ΠR��E}��yg!s�R����8֛wL��ܫT�)�x���M-t�z��L"�|߅xw��WLoX?��� �ΣFБ�Œ����$}�F�:4<�K�����yв�
��:ǳik76�0��80s-�6��g>$�l��S�=֖:4����u��� ����:�ws}��[=�CpD��,$�1��|�����FC`����U��x���*�Z��33IN��#$xD��e8��5(�����"��p9�2T��WV����Ӧ�xl�L�7�C�ٞh88����θ��,���F�u�'}k=A�8Rz�l�#�\�)���i�o�ȩ(,���&R�I}�����
�\\	���3���(�:��[KcOά�⣣1�FFt���X�e��<�Y��V �SҜs�={M��@xx����]췆��u�ͬ�7I�� |u9����`'��So�ɪ�#䪫-�����%r������X��������lذ�Am�B����Bs|�������2��z����n$��F��)��J�6e���do�zB�����a���8`GvvO/���瘣ݝ�Y����?V~�WB���T��?Lt�*�f~����s�
��ݿ%������B����4�'��a�C��A.��7�Fǈ%�.�s��7a�n����T(�����ep<�:]
)?�V=f_���.��ߓՠ[���A���2e��/�?6<�)(
JK����݂�G�_�VG���D��(	"L�K�zS�2�XK��|�``t���𾻸��f(S�"�DKK�\��sK0Sߥ�
p�#(?����C���L���<%�?=���8������1�l�$R���#���а����g�gT�2*�P��Ǹ��$����w��`f��:-���/Dlr����y`�oG����p���#oP��z�'�m�l���I�*?�(�����l�����=�v��g~�
�8��yf�ml���Q������vc~�]Ư�_Q9�s0�(o���o+����i����P|�����}RH���r殆�����1}����$e\l�5ᚁ'""���oj=az3�Ϣ��Х�lmo��Q���2��f�s}����,��˫�Kz��?��F�r,<Z�Z��r�P�3UM��7��'R+��B�+�=���&n�$��չ�0>`X>��u.��*`>y��xdd=Є`t��`��ff2~S��9�1#�R�j0N�>�#ܣ�9v�w���jo��[~_��]�Y�
�ho"�R_�=�t�B F���Jkmϐ���� n����9��a%`m���	��Ds�sÀ�n(�����Z���Jo������|�i�����.ّp
���[4����
fyF�����O*"�U��&��eCnŗ����ʸ�?��e�.�����O��`M��1>~��3�S�ִ�ߨuнc��{S��p-Q�>ܧ�B"Ws2�yg�O6��vLooﲪ�59����ՠ��\q�r������O �FV0���5<-�X	�mt�<o���4!���}�s9h~O�TD�1uu���H����1==> ~���1�U7|��[Kl,gb����x0c����P�U�8���Ye�[`��	}= ����ц
�"8I��s�4dӡ{��a!���C�m�����������Q5zjp������&�>a��%g�{�?��?��$�����A�ȧ��������N����B���S�1�}t��s�K�f��b�פ��{"u�����A5�@ǰr4�� �y�	�1�J�.\��b�T3̒�6��fn_�op�~:U��'#J�[�`:`k�b���58��l�M��BkE9��gN���@6�g��[Z{��
�
�$
4e�6}h�?h=\�_�����ɜ�,S@��
��w׮��!��AWB_���okg�OۧoDD�v(5�{��}~80�����M��� x|����9�Ӿv�C�.���������?���j�ln��P��f�U�8�{6�+�k��j��/Q�O�]�=�����
jI���F2���*��+Dqirr(ܔt|:��ME�����
����?	À��[9�7m�#���`D�⪻?%	<M����b���[�49ٙk�<# �������4�X�K�ʨ���nm�u�>d�VI�P����<=;c�L\�.�ڮ�.���}]�U�*>6���BO�T���qzz�'~�9���Ǻo1�++�8~E�%{�3 ��p���k���EC�xw��y��1�|@n�v������}GF�Yώ�;������F�f%ܳ�oZc�K�爽U�70	��2q,u3ml��!�yzO��h��9����%�
�3{ݧ�������F�uj��M�D�z9��h����#�ST���e�FӖFG���9+Y���4W�K���]�	o�U���������|(����F�@�C���FOϭ<���V�6@�h�_���ʊ�fI�E"�P첊8�����c�b������᡹2Ų����P	I����QX+@K�K��]�{�y��ǔl�A${Z�IH��h]��fg�o�/���|�A#�+�b;���YI��R��;Z!C<���gL�K�JL��T�ۀ�4+�n���8�N���1��i�����`�W!���666���
�J��,.BfH��|U�I��� ?.����^1�F�n̑�]R�LX<39]�҂K$}Z��r��攦�/,,��h�3*Oi�0)%����m������o����s�#~���tJ�`܆��n�茀�.��YH�	���3�~JQ���1������ܜ��&
�r���߿���Z��C��b
�2^Ol��PuH~:���ȳpm7�p���`oV�)/p�>)�p��za��i����Mռ�����
� L�'_�L�%���O�q�F�
xxl(S�NO.l^��ٔ���H6�M`R�G���'J�~�b���*���t.[[\��#��y˱���H�~a!KR�������$-����$^}_OO�Z�@�ۈ{<�̧�k��M���#����<�S�ݫ������D��mj
y��J��*�]?�u������6"�����`4�������2b�~��j�W�$ɋ��Ѱ9�,�OT��Ǐ���SN����d��8q���>>\�h��
]��`���c��	��
��K�9��<+�����hͩ���w�Cs���J"�7�5 T�y�%}���a,:�j:���퀰�����q6BӤ53/wHCt�����醳r�o������Ӡ�i��/+�S+����ƀ�5�&�����!�9�l]�$Dꅡ8�Oz�{a���ړ%N��s��c�+A��*B^��Y���å���־z�7�����'�y�����s��GP��eNE�+�ϛ����i��eP���\�3JLi}n
��v���%V���8�>��$�[�Ӏ�,p�]�N%�54u�	��{cūY��BN."����DktM� '��(��y�����M�hf,�|�ğ�����]��Q&*R*�x)����t5�fU�8/�r�@ؙ9,��L0�s�����gZh8J �?�σ�VB���2��?,?�1�Pr�f�5�n�t��e�#�$��$0�]�v$��b�~RW�\�$�!�ŏ*����m6K�3@�T\Z�����md4r�LP��P��6˯������!��B>{�l9�0bH^l�"�)�L�J'5�����U��N�C��XF�Z���\���%��mN��|��.�)7�F���2--Qc5��LU���%/-�F�g��a�?���ب�	6�K#f�f�{��~K�DkۣRֿ�g;����5W�)���"�Y���rګڍHcu�փ|�Y{x����f(����e��t3���н0��ͭ:�,.XLD�w�u	Y� �t��B-Q�E�R�)�E�.Y$�<hb♽��"�֙�
d�듥��0�0 h0BC�Vb�=��zGrx���s���C�AbM3	a#DNʭr%�D���R�� �a�����;n���lm=V{0_Jd�nG)U���I?�F/э�r�f">�ݧl,NCvҸ���d�¦*�0 ��X�����ӂ/�d���ǖ�˫`c�z5�����;�6�՘�4����1a�Z8��Wd�Ȩr��ց%��������dz�/��Ϡ���"4��&��2 ��H@
4���_�:;(zk���*��Ss�7�o]�7��2�/���,�-�Y�GK��D���G{�2���M��_�c�LTQQ�2�;��_il�|����oE
�6k����r|�u�*�'��[G����>�}�9�d.뱾�Q�cû��'Q�kWEQ����nZ1�W���ۥ�k��jS����o���e�-N����1��}�/�� ��JL�r!I�	\�НP`$���"���M��f�=H�"�da��j�� �{5Nz�2�ŌW�)Ӥ�/[�	�~p�g��?L$�	%�HLCl�~���VU4cdλ�*����߀'�Hָ<�{x�26��`��M�JB:E�C7�?�o�:2��YPZ�r�ٮ���N�o7�?ok(��6��}�8߀&��F:j�	�������9���gV��۩��aw�k�Ix8��S����]����<����F�S����\��X4��H!5i͂7(&�'�u4�ב������ˡ�ؔh;Mjs����j�\ঘ�~��B��{}zvAq�������KI�\�˶��ZW�Jت�rsu�N0i�X�F?5�2_�:�&}�l�U{�F7����.9|��]���y��Q1тW�.w�R	n����M�S"S\9�8zBa�B�{=﷜��@��(�)�z�������/I�3�Q�K���^�j0���M��L���2p�64����c
����?�>?O�h��x�y�[�	�!�ѕ����0�Yq�����V~��=/a�^��o�{>�Si���W���~tc*��:�����DҦ�%�::�;��Pp�)�`��+��b7I!n��p�@]ٲ��5B,�qg�z�.-#��[=`��5Z���
�t�Ei蔧�ݱ�=1�h
emK�(���J���P�E�5�rAH���e_�{cc�
�����G���ȧ��'�U�p���Օ�;׻��6�r�h�=9�vx��/�p@� X]a��
�1i]F(*�eutt�6���O5H��W�Հ��ݰ���&ؽ�6L�#�5�Ą�,����ը�{uB��;���5{]�㥓>��"�H{d��Ig�x��x4�ld\A�(@�X��eam��H�x5�¤� e�37W�<*��4�!u�"����7{�
�2��P �,aT���\}�a�� ����ٍ�Xf�
v[j{��g�����
V��nu�b�;<�T�H>���  �(*Snz���b�V�;պ��f�-uJ)�ksF��s��ʦ$�̪�F�J=�A��I����s�,Ϣ��� ApG6�u��M��9b;�x�G���hq�7�R��`�ǜ� px\\`=�T�[�!Z��
Ec���R������?��3������������2<��)uم�W7��˪Q�.�jW�4[��b��@�0~�*��WN͕���-Fꕠf7�]�w))$�����555��-?7ʈ��s;H��ظǩ�<��{__q�� )�\����cM!�Y���;;;�ɼ��xb{ti��9	o���M���LNO~n�RT̨�Ѳd�,�Blz�@zD��Vn�]�]#
䌌�XRp��ė#O:�� ��#NS<�r;���%�yωe��e�<�_K�`�~G���kNftJ'��-�'���;����0�m^��t��� ^�b���[Gm[j'��3%�7c����w��ӎ��i�^��ƯҌ%4�8Ԍ<�1_&�RWr���*k ��4W ������jg�|>�����f�eQ�&���YA�7q#)ΌA�Æ���b�`���I{.L����c�&O��'�^����\P��_���N#C��I��ɩ	ל5�P	��W�¯�C��u��Ia�a��O*t7�1��ډ#cϨN ��>��G�<��~��m�^A�E���� ����\��()a/��6ms'��9x��APzTUV�#--��������l4�;]�h��i�E΍�8�!Ԅܚ�O[)�?3>�W���ga`N�O1qe��T?(�z�\�]�cl?_j[�����Ǿ�\u'�Gޡ]9��Ւ���e����Ç/J���\�6��vW��'-u:	�q������|�������a�LQ{�bo���3y�U�����2�ݚ
9��4�x�2����C� G���u��IP6#��oSC��TL�h��3�4{�Fg�j�|��d����{�v��!��t�%Z��8]�t�Ct|�#Md/��ɤ�S	�\�	����4#���2{^�M�)���r���kDO�j�V�
ngrϪs���:��1���M����`���&wO�z�o6~��yT(�A���b7v��7H�k�,#��v�W����Ţ�������%�ߒ⸢����?����B�p�� �݇��n�BBh��	��� E �ȭ' �L��F��i��%�{,۴���D�y�H�d��Es4�-X��t^˟!;Z#E@�v�xd�M�w����->�r�������nt��B�">���l���ш����^W}tf��ւ��}�2�<(/DOOO׌��-�g^fQ��'yj�W��[f"M�!w�&|ʲ*���%8����s:d���3ɿֳC����G�g���ҭA鏉�kLa���o���e5����3�3+7T=WW'HJAB��M�/�U��gi7l��.���eWԔ�5�g9���Z��KmU�vǜ�X�}C'���C��¯Ǎ �#wn��eH�1'?���������{�ۓYߴ�4j:�����O���q,tZ���7ϥ�Rۢ9��o��~��u �/��}�$�م���Q���B�����]�F�P���q9����L݆�F�u�o/��-D�;� ����2��{RT��Bb{-u�(�����W��--¢�+�N����LG���^s7A� ==��G��;"�D��x�Kbrj�j�=���?Җ � '��33W'���&����hD��8oJ|�XR��8�;)/�ۨ��2��Et'���L�,w�ڍ�z���i����}�N�G +��[a�}�T� ��0��n�n�p/�@l��ܭ�mT���:�R�Lk��B�+������1�w:��`l��������p(���2E�9$���N.|U��Go�
=.���GI<a3�����NNM��ބ�����y
��t��EAw�r��턖�B�+�)���]nK���SE�`��̓�Е�e�O���ds!��J��Ô��wt��6����G���J2��E7��׬a�/ŀ7���wI�V�JiNƧgكP0�k!��nY,&���.��t��2�
��&��LW@��:��+� /n^��k�`"B�����'�`'��~R
��D��I�����0�蝊�9=��Z���� 8�>*�?�Am��GJ+����mNw�H�W�^k�����qδ�ڒE�ϽW��H�ݷ���oD*��A�P�3i�@`�>�k$x�)�@tHx�����ܢ�(X�^�ٮ����FB�$����������&s�3wk����4�����}U�b��L݅�A#��дx(��O����L3�F<�zO�2J@����Z���46Rmy�S[�([B(^�ܘ�[��~id[�ե�y��t�]Y���en��R����� ₙ4�˪��Շ�AJΒ��!��3k�n�G	}�U�p�ʹ�����1�P��� -�K���K��#�jg{i)�kF��4<L*Z��cY�������.Z:�N����B�K��s�[�&S>��y�-������
�	��j��@7�CC�G@�Ȏ��TT ���oBZt?�[W���G�5��f���N��8e��?��D�X�.�<���Y�e��9w����<���6X,�˗���H�73��E���XILiZ��p��k���j��6g��/eυR�j�!tN��Rܙ?7<�/z]�zg���a��90�V KJ�fi�qz�c�H0|ap`�)7w��w�A�+������M��cFv�W�Fv_(�}KH��ܬ��5�k��a����z��@p��v|=�ܡ`��9#V�DܠUk0<d")�=l)W�)�?�M�z��j�y1��j5B*��խ3����ak�n���X_�P�nOX���պH��w�g������d�9|��� ���r]�����`[�������;�����J�H��q���1���}��m]����'��Az�E(-h�<,xou(=B^���)T旋G���f{ʑP���X B�~2� �k<��ק�G�m4�
�L� +6�D&����V�>vө_�O�ܷF�!yo8�<d�>O8�O�`�����W�
?�����`���%Fm�+.nΏ�`[u�Nq� ,?Y��~?����������D�q���>�����y���q����+թ���W��/[����:�k@�/�&�<�N>�I�qrd����{���ɳ��\dF{��'���9�}�8�I] 0��߹L�V��ץ���I�ȏ�	��l���� ���E���c��B�(ˡ����]��n��*��`pj[���ʐ�5#ml�+�¥�U��p���0�zAq�P{W�d�����4��������ꢚ��녙����s�OqTA���E1�c�}���E��W-�䵮o�k̉�"�PJt�K;�㛪�y|�������P�������R������ ��e/���&:�н"5]m���A��#K����l�`Vcީ�+���g�U�h��p`�������f��6�yG{��މ���M��B�>����f{~9ݳ��-�:#;�cI8�A��ԙ��0p�� W]�qJ����D�Bh͔OSKb$щ=UW�GV��N�Hk��6��x�"�z�W$G؞��ވ�WM!�5/(]3�}���x�:���0:��-����/o�K'V���q�&�����?��$�9�^�(7����yR��*�X�k},N6�#u��Ì��b"��8�����U����px�j���?*'�OuvJ5�z
`�G='��I�7w!�D�L�߿�GmV����9�eq�8�� �ۻ�W���-�r�����fo{l��||ITf�?�ٿ�!6�ب��Eh8��6F��<էi��V�4�����^X0�tSѫEU7�٤2K7��T����－ >��qst�p��Xg��f�5*�A	/��&0���pky�t�B݊�?	9�6�j@��26;���ȝp;!$�L���W�w3NqS����?�[��Ү��٦Dr̘�ɝK�m���B�+�R��X�����wU>�454)���Q8���&�˻Y'%���54
u��`�v���@a�)�2k�T��/���&TѠ���������a3r/nD�6��ѩ)�����*f�N��R�Tu�<t�i-��dV�B[�����y#����9�}4�`��#%��DϜ{���.�M-+fK��%w�0Z�:�RQ��<�K0={��&Xz��`��$�̤�� 7�Uw�9�.�T!�=$�F��A*�?��uߐՇ2�����K!$r��O��+�1ON��P8w����"��#x����2��1��Ӧ����kd
*����t0���`Jo�g� "M9R�Fm��rY5᪏�%�,�Һ;S]��]$�/�hl���R��ƃ�53�~5U렌���S�Ijj*ħ&��̓uV�}���9�*�:���1�����xb~��ܦ�I������9�N������I�����؟�_q7lo;O8��2��wp �E)P���]�72�y�{�ݵ\Q&��uL�3k��3��444�����䕞=�	*"���S���61j�ƅkacC�>�w��,�?�sȮw��0ͬ���П����]t�$���E<9VuT�}�n��d�3���{B���5�d]	�%S��X�'�N�4���z�ڕz��w�Պ����8���p ��z�И�`���rp,����Tc���ǀz	�3�2��d���갨��}�K�����N	i	�KD�N	Ez�D�F@��a�p����}���~���R朳��k�u�k�䞹H�u8�=P�k�؝m]�AX~�l�����h��� ��|�ޑ�PRR�e'\f+�6 ȕ0�?�0����oyg�-$�o~⟜������P�,�������㣢�9^%kG ��� �$���P���Qr�[R���S�C$��Zo����ֆ\n~�CU��"��qx�F��:�h%��x\Q830p��C~�A��,�<����!�X'�-�O�c?t�bFΗCr�A�n���t��0�lb�`R����s���f�l�g��{���ΜMнeȭ�;̬ �Q(���������0D�`�8�v��a��ʜ�ޜ���Q����P&%�u.�Ë�ꤊUV^���_��X��l�����D}Zu�U|���igZ���j��M�'AڝתS�&�l��޹�����S�������ڵ$�Z�_m͗�_V-
�P�K|�v� ��QD�*~z�4�Y��7Jː��8���R.�|]T_��v�EssV�z[��W"��dߌ�9͉�(� ��/�m�[1�(}v�72>�=��I�@��~���ҕ|H{���J�RFv�i�Ϝsi^�͛^��D9=���w���`�QH��Պ��(O%PVV�Ȗ�`�� \J�r��9��Y���D��z��P�O������kxe�44��F7������/I���!��-���a�S�R�Bn>�=x��e��&�P3�X�������V�RG3����!rK�+A���Nk�Т��L�X;�Xcˠԯ������f?�kf%�i�躅u䴢���
I��Z�%ߍ`���s�R��]㺯t�_L�e�n�^��kU}�JK�^��$@�u���3�<���Í-����Yվ�Z������C���p6n�`X�:�l����Z�?g��+B�l?%*Re{���o������Es�N�ݭ�S��㟏u>��uB��'4(_��Ƥ$�+�䇋"�g���p	�^���S��|q:�yό�qe�����rN�iӐc�f�ڎ1Vp����M�`�A��ϩ��o?���`��_$�ГK�7�h�g�]h�Z����q]ⲯ��5�vB��0XR��z.'H�I��������5`���r�ҟV�`��Yd�;{a����u����:�Ӷ *:�c�l�	�$X�xh�`Xa�B��r��$;����E*�H�B0t��Uݪ��3�&ަ�9�5)V�h�f�;_y��fyD��xo72$��i��;%b� R���16��D�<� ��\ol�5?���N��+�S�(�B��>=6}�lᡱ�����E�%�hVxBQIN�7���JN���;TAS���E��<��N҉O�m*�Չ�FЄ!���Q�f�����CC	N*e**0�$�E�t�Lh�o]�_f;_O@�>�0.��5�;;�|�����#`T�͉���*J�ߛcN���D}�L��q�0BGd���� .��?�Q4��\�>��2�9)76~�V��݃��
��ygԾ����0o-H�6b�(�M��돧W�N�Po0z�Ɨh����������B�i� ��� �$ ����Gf�	��<����L�dt"���p�r\ӣ�������q���Q����,ǽ�T�H)4��6yz��s��0
�`�PQh%�k� |�1�Q�fX V���g�2���ǟ�	wkk����Z��/��1`�qgЎ��زO�?�ߝ���FBOF�0��U&&<'UERM �鉧�s��q�ݢg�C0u���0����-@Я��L8��rڃ�/��V!!��{�BO�Sz����� w(���U ɩ�&L�]�]��˜�Y�'�� n@?W�lӋ{"����"ĦE��������&�iǮ���
�Z/���`7��wߖk�++{���)�]�o�;�%�`3Jc�9�o�)�D9��J��q3W��ʝ&���M0�?>~�7wJ�em��IS����'5�Q�/K��/�?5�s�x��5dvC�>X�X<D*�*Vغ�}���K+w��o�����ඤ�u%�c���(jJ�CO23�q��tji���E����0��̎���\_T���e~�n��q����\[�Ą86�f
Wey�Py!^�Q�U��z�~pM�O_��ݣ�!���F]�C'?���˿U�8	�|>��PO�c�@:%a�gT���{m�/G��_�jJ&PY�_k��s��
�U������9�`�X4b��QqQ�`_vu�L:G��7c��-��t��z�5�h`` Pv^�o���M�t�K��#�&������q�07+�7�5!���ؘ4�"%��)`�%<�~��'���wPx����������X�6ii�F��9���?�^#���U܃���ma���_L�..*���4������a��yp�-:Ue�Cp$[,��n��Uߠ���`�Xի�����v�j�S�� ���>5a��������y	�v)Ʀ���HȮ��V����������{�-��k���.�2˘R~��	��ލ��U2��Q->	NNd�-k�{�QP���3�}�V��C�m6L I!Sssv�|^�h��%�RǇ(��=G��$+�%�W�p�К�P�.���@�W4�q�}p�'��.�G�w���� �%�Qŧ/�(���NN5�jtwen��ek�Pnn"��<�ed^��Q�d"l�m%�2H�(^�x�p��r:e�C�����܀��:��i��"b��K�|o����j]NZ"5şf���o����sq���",7Řn�f>�Le;]ͦ�f�f��N%t�!�i����橈\��q�a�'����D���q�(��>���|s;�C�		`�~���[�$�Ĺ��d,�>�W��mm�!�o ����=$lj��1,G驎�f���Gln���=���C#�WM�؇���X�Բ�֧�<:WU%YO)<�&`׎�{O?|��'�=bKR�0�I9�~��]��S^�D^6�H������o(�<�𦢭�⩧֭�q����\�|����jyL�P��|�	}�_G[Ӫ*�?�/��]��Ic�V������e��a���a�S���/m	z�'�(�73s.W[\��f0���ü�<<(_���"-�	��4�A=iL���0$t�����*������rsoL�+�T�87��r�ZD�R,ĒΣ٨ölg����4ߛ�,�ҿ��@j�Y�C���$��$A�{���vu>����9��a˄h왚��t�\]�v�p���/��@�S��K��NNOc���M��%�2��S�Vx!)UT�
6�D�*ۿ�եt��(�(	���^�Qo4���4��PW)�:5e��z{��(qV[�KJ�A�ŴEp���S�(�_��nn�.O�;{�ד���P0Z�+>���݂��l8~S��'�B��d$�?���(��J����v�nDN�yG��e�mdX�Fe�\gY}tN81�;�Ã�3YjV���w>ĝ��j)� �4�Wz[e��C.�刍P�j\.�-M��L�x�k����QN���/�»WǶE��^(`�u�MXm��cb�bŤb��uZ��%r�v���.��9jx5�s�K_f��e���u�;�*A�E����سP���<3��2���sǴ1m���s�$\QQQ�<T�FB��D�$t���r�C٫����p1]���3��C�,WK�d����AX�np��c8�?dz���2��?�K�]t[,J=!������\�̔��ף�K=sS�'v�\���,"|�L�*}�1�Vd��� �B%��Aj�3�6���c�/|8;�V�~��b�n�^�	7� �#���gY����%�@Օ�Ƨe(�j�N�����3�8�Ӝ?}�S�6XGK+��	P��(�|p�?y����:���!r���ug��W�9�ў�ڝ�#��>;;:��
 �O�H����[��������o����$��c-�UL�cr�v�V ˉ��2M�FL٤t������KZڦ�X�&z���ͻ�[��-b�I�,4�ZOǑy/G��!�A�;�-m$��� ���z�dif��O51/�*t� N�U|��)�[>�U�e9�����d,FOf\��8|	p�LeH���X��#��6��y�6n�P�5�x0����qr􎎌|((`-�g���TbS%�=�]h↞䮁8Q���VZ�������� G ���Et�34�fj(���#ӆXg`|^��Eᖦ��ˡ�Д��{2y�_W��>��!_���\�8F;l����>��+.N�e��k�y�p6���e���,�r<��G<{���I��	Dđ8�|~��Tcb�1@4;�����(�a?� �ˍ���#���Iݟ�Q>�K$⸇�����IZx�.�;��� ����U��W@7<�������U"��l�[�X��� haV�@_*�J�Ad��m\��b�
t��r�>�Ux�]ז��ɿd�Xl�JK-`>�����F ����Y>^
��`w�i6),�//����5i�K3RG!ϗ�B�$짮��u�6ԩ#��>=�H�'�Rt�z�In*���t��	8�km�Aލ�oս����,>��=d�~@�;<�&���&�@�Bd�w��n6�x���܃ 4�K;�R3M�N��`S�N �?���0*�K�[��%s�xy�B��Zu�����9����)Ő�ғV>]�>G�l�����&(��)���$�Z��+C�1~=A�=�IkE�pg�f3QYy��0I��+0ٖp��C��I�����с�ֵ���5p��š/_b���i�0��E�PU��/�K�\m9�s��� ;��&}�G�1���~����|c^��]S/���<q�&S�24V?�2R�kiky�-�>��A���B���$����,���|������lx���<�0�Jy)u+�	zN��L�~�<Z ����<��D*�+�=��#����6��=rD(ڟ"]��U�@���e}���M4�� zb����Znz��G��x��f�(����ic�r���K�}z=�j�zl����֒��⳰l��T�i'�Ѻ�'s��~���C@ƨ�_`�l����q	�U� 鎔��(���l�I�/mr�|.`�YK�T�!ς_*�1l���`�G��O�_(�)��LN'/�L��"�{��@��9�'v��(ד6A�L2����Q��y��8��Ҡ�9sk~~����e��	�5��QJ8.n��B37�ㄊ/<��?S%,�#���+�=L�b9e�׶Ks����%�u��j�-u㊉W��2WWMt�x>7~_Q��jk�~.�bc�rW��qib;�s�u�H�q�g "�p<6v(/��g���8ͫ�m�އ�2��m:��d�:c̾��}}�����"����]�/������.�O[�����q��Z��E�*���v��RI��4�	��1C	��n�oK��Aa`ϛ�u��l������}8�B�͍o�DG�x���/'���Q>䂽x!�s����l��xZ���E�T�%Uo�k� /��L�y�0|�õ�ɑ�@�����g	��u�m���v��^{ҹ
�/��Jp؂�/Vο�B�t�1^^��_�Ix7{���~l��V|��s��H�����Uê���.�J�Ԥ���.��#QGo�̩��u`���[��]1�D��g㓞�������s�CT��D����M�;��L �2�D�o&o�ؖG#���n��>9[���A������e�ģNx��wy�%�� 2p��0�Sa��!mĊ�=ih軕c-B{��$�v:mI}��楖��Z��[h�M��a�i�m�.r]}�3Ȝ���h�<	3�X]0��`���w�fh�j�x$n��Јp�7{7�c(�w�_����25����������L>_X�3z�C�*{l��(pnO�9�'�W����]�q����!xrϮ����{�I��X�䖸����m�$۪CU�N��*s l��2N3�h�d����d���O#*z����El�7�z�[����JC�u�,��~+m�e�'m5�>X!l�|��b=$���_������gh$�K���N���t�ޯE����*�Jͧ0�Ġ:ҿ��]Q$������[�VA�淐�E�+b�I��9c��:Hv�'Q�Q�S�#*V�j������������p��.W����"��W�GKP��3�G%���gS�ќ�
%��h|9Ei�-*�{)@q�啪��n:�H:b�Eۿ��]%��kf���Cߚ�cHz3��j�\IIi��&���l�?xo]Zز��-��i�����YϮ]&��EsoZ<�����U��µ{�Hw���wkWrq��r)u�-P�����L���;�H>@�����Uj��S�[�/o�kwE���D�RG(�����s��nby�59"�WW8r|�`�}liR�G���"�|��˿���Nw��������sȐ��率㼏+����>.�|����#�U���l��֐���c[d�ͣ���>t/G#���+�����<XLy�P+���_r3/��>[�@Ս�V�FY�&]>mdU0�V��������u��Ryί�D�b���lz1�OD�f�#33zzT���旕9���2<?�.�����j8�a����,0� ��;����+
f�ީWs����z"S�	����^u���	�7X��S���zqPҵ���"+�<�p�ۇ<} �ʝ�%M��/���x��̂OoEZ·������um�����b���0����o��B�ϗ�ۨ����Y��{��⤱|�5�1i�㮫c9[˿?��}}��!e��cZ����h>�H�����i�A�"�5�1RM�����ї���&�88�%�W����\�0J��d�7f<m�&x������!���#v~�SӊvJ~zw���f����#v�_8V��*���0y����v��c��w"��C��˛z~3	���c�GG��b�z0�:U��}�_ ��^�z����JhM��2q�$cA�����G�:��Mpp�>{���y|�wq@ꫮ��{3M�����'�m��S���5���e�)@�`R2���(���Q�➍W�����^����N�
�f4�_!�!�i(�Y����g�Ow�������2n}��W}"��z���m�[6U�V�e��̩+h�S]��~�4� ��Ub�p�)0�G%f)����2<��WL��H��%;lX�ތ�������oE���E��Q,��I���7�?v�NX��(p��Tm)��!g������;�6��$������_�	�Nr���dA�F=��w2�F�
��,N�0c��c��h�pmӷa�B�25e1�y96F^RZ�L����?L����K��zaZ�I}�f(����x��lex���?���Ⱔ�c�Z��$�5�0�c*-&��0*�^^..�g�&�Z�H������`⢢�ã}�@��(uc>�\p����kZ�H�NH�rpp�0A۪=�/d�;Wt@'��X�h&lq�;�}~r6v�2�yV�/j�p����M�!�Ñ�
gtz�rD|ir2������ �=7"b"�[Ծ�!{B1��GNF�TA��];�N��PM{{ڠĶp���O�Ԭ���1���������� $sH�vC `�W����?���	Ί7X�_L9��u_�X'|1e{��$>�À����W�1����"���?�\�3f�/�щt� S����b��f�4�j�J�_p�|�[w�.'�,�
c�;l�A���K�������u�d_�7W+.1�0�,փ�A�Vŗ壡�yA�����pz�U]FvZ��A`�c }���uޞ-�V�T'���~��
E�W�F��6]f������5��j�_-o�T@��K�޿�z:ͯL��!�^�'���@��0�c��Ą��T6��0+6r�S-M8P/�����[w�{�z;����ӳ@oE�߶ieM��K�����$�=0P��W3?7�+�T��O�E�_�Qz��S�=�+��Q���u�6�,Wa��s�z�|��[����� �O ���@'��[
P��C8��p�s&+g*g~?-��q�p���Iz6�,�Ͱ��l��[ ���C�������'��k����ֱ�7r|�8�(0,�ZRo_{&)1�h0�jJN�����p�C�#(.EO0�c��K�Zt���������z�ٜ��ly��Y��W7�1���Ûأ���5�!���<�윤 ��)W~�Z�98;�<9�p��6�H4\)���&ATgPw��L���G� H6Q��~�%l�"qS>@�QWo9yڐ_^^�8�W�Ho+� /W�/��,8��qJe�^aF5�gg�����P$T	����a�iN�����F�HG�k�}��&7�fZ�KH?8��%���mv�����x	\-nOLL)��{�+��6J�q���3�cn{�k�Q��a�$�C��#�4/�pTs����U��!].
Z;*�ȕ@//,J��d�q0��6h2ɿ�~z���}6pD��=��m=q���E�����{��jGV`����a�A����@�Q�9�U/eA��A��H��!�������d�p�R�?� ����.A�8߳�PVU���LA媴�@2M�W\���
0<���O�l����AbجQ�~
Պ}C�,�kj��OY�mS̛��]<&x6��h�k̀K�@�9�j$G*h��J擁D��K^�ݴ$(���'��qX~h��W��2���9��U��� �}nQ���.��O
�]�~U;�#pC�qw�y��R�TQ�����sW��	)����ƴR^?=q���-���h��un"/��>�g�A�����4DG㜐���"�I��t�nr'v��*)���M���w��S� ���~,D��A��?X:�iM)�tb⒮�N�݆-~C���㪢��dKv��6C v�Fq��
s02{�l����V��]�I�46�6�_䐸���Օ�w7�E`gw�#غ@�xⲲ�Up���ʆ����17����Σ�>���&��W��N~H{�3�y��;>��W��xե Ҕn�REL,��ŭ�Zo�c���Ÿjjj�֠wA���}���ۊ?��/�y�Y�ےr����\�˽�������<|�D-PrXD�5#�(��،u�n�G5S*E���2��o���N��88:�q�8�	��v]Y��_W�Hmb��� �b� ��:o&h,~ײ<R�@e<�\L���yN�m�F4���\�<Kћ5Yä��k�,ө�P�)}˗/���O��*�.�I�_�ւ1Ҟ��4����~���"III�r>d.�Y_+�ǋV�a�S2|/���寡�7����dI���+�י�5�:�.Z�s�#3?[���&\l~۳�����|?h�w��H�,!��zh���gU����	DxGU(���!�[@Q�������t�ê��-j�#�~@͝0�3�Sߙ˼�;��I�b�"��E�pЮK�yo�7�x6����q��c+�R�����ćƀ���ݍ!�"� �NMՑUɍ��{�`�ƣ�x�ׯ�����g�����/o�t�UT��n����嘺����(�>1�Nm=m���BY���&���F����Rا�G�̚·@�:P;d�K�
�4]QRb�J�E$2�Sx����q��[���.���wxa��#)�B���`�5=����v�F��)�J�Gb/Nx5}��|���%��@�*��f.��I����h5��.P����!0�tt�V�\����!Z��� F�?�u��g����|�ؽ@{�ƚڥz��� o,���l@��,�%AS���Rh����aO5�*��+yYP��Է�H���>;���!�2�X����[}Z��,+2����q^Y�~9E��ʏ���X)�3�U���ц�+4�b�x�L�h�sQr�Z�c��� �u�YYY٫)��_Tid]���_��I�	�1)Sgj�ِ����Ժ	���K�
�|͋"6 P�U����0^�^yU��E:j�bo�����j��(轥��nƚ���<�ա�j���";{P�ؚ� ��4�:��O=wvº����<X;�MS��o]A}{l!VC&���Y7X;�+�yDb"�H�G��&]��R�t�I	���8�ƛ�����2���'Г�p煚G�ax��&a��Ѽ���OZ�xDc�c�ߑ�ӕr<~�^c2��nT>O�<�f����/����H��U[q��qЬզA�0������K�y�6*N;���J逪d�����ݎc��W���#��]�{�6��eoF��J�vd�ԁw��kZB>Vw��r�j����&��'F3�v�4����2�`��'L�*`Q�7ب�zj�����zoJ�~��?��[���؏��Oߟ�JC�О���"�E�h��V	�	@�^����dhnn��P�����L����������n1��A�'i�<-m�Ia}1%!!���)}�����Y�g��v�����U ;9>��\.0�M5�L�A<��{���{���� |���v�Ys �%j"#��.NC�A���ysa���O��h��h�!1dL��"C�'�^�^_~z��щ��WZ������������u�;���jL��q_ 6�|
# �Ʒ%P�\wчm׉-3�f�>:���O�\8C���깙P`�ғ��ړ@j}��Jc�|Zx��9�&����Â�%�2���9$QQQx8���d���L	������������T��z�������C���(��?��l��]>�p���q/��Ģr��#Jd�srr�%����LX;�i�N]Ö�3M����~����Ⱥ� ��$o�+~� �xU��M����e�1�P�n��ػ�#t�AO�B$�Ú�J��k#T��J&E���*��F�7�����^Dr���� ��[�2���}tt4�\��F�v��(οݠ@�`bU[�����?��spr��.��ÎP�\�ᛵ>��fn/������&�8P��F�����_i���ج,Z�y~������u^���M��-�c�?M��6�[Ҍ�%�wO���o����b����a�8N��Ae�h��ZS�)�����9���JJ���X�ڶe��¼�P�C:�*��H�$UE+����n�#�9����4#���<,�#S�㙷Cξ �d9�y�����?���g�GvO���*���aq��<[%�8��x�lR��2��$7"pq��G�뚐_[!|^9��|��5����X����ܜ��*P��v����Y��f�� v([&J�+�����xe���m���K�Qb�����K�ʿ���%�xF[m�I=C�=��ȴ��7��};�N� S�)h����P�t����l��u�{Y���B���T��ϯ�e��'�ٙ���k}�w��7�G�@�]�r��m Z���~��h�T��9��ג�m٨������a�$&�{�s!��N<�y�߱wޖMZ<p��΂E���&��֒�E���H���<�ΈM�6!9A]f���3+�
�6�Iw������Ǣ����#������]��N�E��dy���=Pm��u�ћ����8c#��n.�1�O:�]W���4�Dt2�~{�^f��67�t���h��!��n�;�]�9vUTXy7;���͛ 耵-�C"e�67W,UM�	�hݯ_����,;���LU�4�>۬����1���LԶ�ekp��jU�6�`� ����rC��+�`
fi
�fbQ:w|�pٵM:v����DPL����������b�rc�>4����W�=���|���-�y�( #vv�V�p�lI�=������ ���Vj|E�^>�1��Y��Ve'��>���_/X f�b�p�I�pz'I ͂Y��m�)�n|z
<�/�R��*Y�}tj��;��@�R�-89ڸ�����	+��Ӧ��0>&$�W�O�����r]xt��'�7���`��ae�N�ڥl<3�^�׉Ɩ�qӟ���3�Pi�V�_aQ�hPZ_��ކ�W��Ӻ���DH�+e����_��ۋe�O?�t�7)n�#�&tHF�F��Q����̋���>|�}9���Y_��q0�����B�!���Iʖ�e��կV�V����7=�_bB^c�Toy�b���2��24|�.�/YS�`��X-^��^�$��9��nkT@冧��~9��������� ��	����<��v�M�MMM��_�����G���f���c�H���T��\t������	�����ď��?�	�B�����(��=Y'|+��$Y���^$HAH Ld���e��,00T<�2����#��������#@�x#8�<��������ρ�F>���"!vB^��c���q���,��?��fN�~�Bu�$�5��-�[�~(��Kj*�� 5�7o¡'���4:rH"����;]�T,�����3�f.{����	\�Il��JK�/������k>�O8�����K��srr:�̾~g'�߉ǈI̳*�=?۟�S�u�@��\�o�Փ� 3�t@.:�B���^&�)�.8��ߓ�{��}���<����\w��s3g{�F�K��������i�W���f���g��O�
���4�0t)�y�y잩}��A�k�e�-����2��Y��Z��[������@�]G���\��Sy����",���R+��Յ�ӵ�z:�z�V(�����nu�"���_Def�P�?|��I�V�٧��9_Wm|����ǷV�r0��M��u�{���̀S����W,`�e�:}* ���4Q=*���A������M�_�i��'E����~�K ����P�G'��G�__�%�Q���|� z�G��5��ҙB��jB��z����p��|��&� X�S)��R{����5��>,:�����W�O�w�����ס��#p�|nn~����K ᇚ��LagGť5*4Ƣ슊��sz��m?:<WU)�M�Mڶz��]�:I����؜'���"{]�:IH/lhHD9׀��| 	m?�N�n�����Q�/m�H����d2^n�g�w ��/D<�90b��$�ݿL\����z-���QШs�9�'��N��&��d5�d�	.->�TM�O�I�;����Wwsqa�:!{��H���[��h���hhi�>�'Z�[�풋��"C9�mťnk�7�y���a�c��U2#Uʇ'�|9��Sڱ�G/I�j�Y�"y���+
@���Y1��tK��]���SR�m8��֌e�8K�|����'p���}��h�!g���s�N�L�jr|?P��CƼ8|s�184D�?��Xb�jH뭻;��١�e�^������ƣ�0�?|"ö��8��Pk�E>�t?�xXd(碳�R�$3y��N��HD��M�L�]XX�{��6��ށOà�{�:��rk���������dk '��wD[�#V��E:4����'XI2ﲞ	�b�(�m����5!V�d^��NԨ,E�����w2D�%�ˋBG�b���W9�-���׼�Dz�z�}'�;(PXV̡�K3���K0���֖�wjLOz����"�A�k�nm���%��e q}ٿ��<�q�̽�@�U�����tK���>��`�C(t�a-����ش�}�-4�bv.�<�Âe��Jx�ZQ2� 9+k��!�*�����uVV���ݾ�q6.���Ir��lq�����?(��:��z<e�k�H��@�����x�.+)�+z�2���ǳ�*Ӿ�lC<ܢI��t���IǺ�:V
"��3�'eq�gB�䪖��Y������"�z[��N��K�N �[���<��s�{j��՝����F(8����G�
�4�ž��>���w���3������H�eJ�>�~�]�ˊ���hR�韆�HbZ�\���j�����" 	�y[�SS��)�*T
h�_\eVl�(�:��D�l�Jj�?�/���F_(_��p�M�E�YX>�am��U��2�?�O@�ؾv^p?Ӟ�Y���eJ�
���N�e��[��J2-��"{$�MQz5�u���>5�훛u��N;�t���[H��`�a9��X*�T�)i�i(!��c��A��\�@�H�����fuɥx�%�=��I�(ҭn��6�=��aN� ��k���ߵ���6��7��)j�115M��歶T�3�yey^-�r�'L`��1o�����I/tf#�B�]�����埝;?8���_p%,͆�Ga5�>��H9(�Y��ubSUx�l.��>�y�w+W (%�Ykʑ�H`|�Op�/	x�W�2i��o�U�nP�ݪ��5:�E�/�d'&'��j8��HM����W�Ρ���%��9'QQ��L�vA�!��/!2<f�$0����z6����*z�se6�KA�x�5� ��ޓR�G,5K��S��������N1��Cj�88B��4K���;,���{phPHj�1	�$����G��`m97�"\L��Go��U��+��Ds@��Bݗ�l�q������LX��N���00�D(S��R�6E[�B�"J���vȞڠ|v��������a�WÊ�IG����:�B�<�7*sP<<<<��ƪ�Kf�&E/)��D#4�A�A���;��8�7�l��@��d�U%����O	��.ܮCE�,*Z�i��>��#j����hxPS����*W���.ܥ��� �� Z��?����a�3z�_m���M�؇l�q߈�� m$�9�E/�����آL�3������7�ZrqQ^������Xi\�(rR#jfZ��8N4@J�$1Z-H�	�C���-[���G�-�B�����.ܵUY?u ���d��O �{�P�97�gX��%���o�nT�����Q�N��ۓ�����W�zF��$TtZ��Y ��.bHHH(�~�"ڕ���Y��iA3���Ś��4��������..O�=! L�}�ݛ�Pl^�?U���i(«��eFvNT�]�v�0��Z����<'��n��3�����D���1Ў�H��֛���&��A��<�����a�����hk����'�Km����	=y���I�D���Q���c�Ɓ���}�^o��Ua�+e�Ȭ�k+5kFi�\�ڈ��& ��7�6p\�g��˹�#%!��Z@���2�%թ��M|1��)��9�A	s~	����B�ԑ3[7��0H漣m�p2��.��������\o�ᇐ~h�!�4߲,>ާ͈�Л����kzF(�^�%i�ĄI=����daI}z�is�[�V�(\V���i��e��4c�mp0�?�e!R�o�h��1�K,���n��*�`I�X��(�ϖd�r�ӗ@L��B������^���;R��Ь�]�0͏}��
3rr��d��|Y������`T������ogL��	�l5����|���$.u�N\đ�)V�v������¨C$f������ 0�b��)'G����}�DnvvD��<;���< @(��	��9Y�����""�Αht�$���]�Yy{�HV&"@��֘Р�'~E�\+X�@�}M���7s�C�*��n�X�$�1(�a3{K������f�d�i�� �>�y�������#"�K��x��Yi0x��T����$Yr`�µ��~��l�@'���"��<�<����2�m��gr7n�Y?��op�]�}fj�2rR�Q�����/S�UV��#��Q|Rs���aN_{u���￉�԰[��C^�UfH��aix�A�r�|ҷ������g����%$�m����9ܱ($~��΂J�q
�%K���甘����\t������r$ܚ0.�'���`��]o荡��1<�(|bR���2o]�9`��Y9{���E�����တL,	`X�m/��w2~`�����e+~��/�nڵ�OM��������v����>�2�����ng/4�O5 �4(z?�P�?��Y�*�PE� d���I���gQ/��o�hX:?'�t;�#�,\����\���@�W>1h/����)��w\G�;`ѵ���"�r�`�he��U氌5��+�D6?`0gŰ�m�y�B��6]���@�03�0}�Vl�%%��2��0F[Tǘ>r�A���K�K�,(%�����5��k���������kc됳b=�8O���^��M�Yav����?6t/�����hbZ�D@Գ z�/ii6=q�� �},��e
�ZiѮ��K�/O�\��om�a<.6t���>�?���Y�a�+lgˀ�H�ʧ\���m����&�R!�q]����Ժd�ov>���3Ɗ����`��%�����穻z�z�6��
EQ,��k|,N��z�*p�kz}s#��J!����	��n/��_rڄ��|	"V�.!�������jo�t$�+o�ud{vD+2�~��Qp��_�ua;ԛм�m��q�Opprz��8���2�#�s&��f����`ٙ�s�=��.����́[�D���c�$8���]P98_�Y��6p��50`��Z�@EE�̓%Մ��������������a>a��G�H�!�����W��B�j����G����t�����V�#I%%^���:6�r~v�.�=�_�� Ю��m�N��	 ����cbb
�gbb�U�r'��O�D���%���N��?�:d�ߚP��~��<�4y�M�������N�>H�w��7��H?�9���A��Ҵ�{k�ɽ���vpЊn����u�v\��8.h�6����;u����;���òL(`h����(������?�a�������7�n��i=��x�23�!���twzdlN�4��LLL�p�R`��WOǟߝ1`� �gdea$G#�\�9�0Iy	5A�瞦�.-%r�S �(Oc��&���8�O+M��K���G�[D�E��twH)-!�-�tw( ��twH"C��tw���!��P����9�s�G��;�^�w��bVv<I�q�ӭoӃC��GLf]�$��ƶ��MC!�ƞ%p�2��lOVؕ�����WA�<��ޫhf&@�X�m��,@T�j����(t���̎�V�|��fFe||�2�E Z�I���G(�ʋ˾���&V�������;.��Uף�j���� �𠡾߉�>l�a&3��@��v iq����F���糀�����7�i�f�I�O��\�����*=1>��k����;�!�n��h�g����eD..�t\m�m�@ׂ�Y�d�Q�tO��q�?�ziY���/%I���V[:��" �f���)sKWnP�q_
$��.�:��Uv���a�HN��Xq��O1RG�����*�j������g�z�Y��9&�Q��-��k�#�vD6u�|<���L�'T��{��1�B�K�"�q�{屳,r�~¦�����G�$�@u�b�7��DK����"辻e�q4K������C��F�@ Ey�K+�&�4���u��%d��	�6�� ���"�q|��QJ�{t<�SsԊc���N�&�p��M:99j�_e�=��_Z��rF�΁�na<�ee ����m/?��O�IN�z?��-RU38��#�z�]�-�U~2�.A1Ņ���p��`L����߄���FQa���
����$�����sA%2c��4���Z\�9���p��'��9�*V�XoDCZ��0�E��r�q�kk�P�&�����P�����J�r��4|�m��Uض���7�̃�Y9��:>��͛7�W��$�d��C�F��\5b��a>����1L'����,������
����{V
��L��G}W���O%%	��5�EN�����x��"���=�9��|�v���m�~��!�^l/�K|�4�=�7���=��\`�Pz��)b�>�-�Re�\ٹ��������<B�K?M�aSE���zmj���6�G���}��rG;ƽ����eԼ�T�d��2��ؗ\=4;Ĵ��ס<Euc�|���`>�S%	H`>�r�k^!w�Ŀ��<�5&�ߨ�������X�+���)d�������O:�9N�,����eű���V̋fW%�y��}T�ZZڍ��$�>��w��(0�DE�o����fg*5�b̰P4mT;-�1b�gϞ��ￖ�MVK���#�T���²��uIDi�y��_K���!�dE��l�
M�IL+��-�H�����i,���WR�u+X�k��>������;*� �0@wl!��Qw����5Z�)D`l,�b��j\a��_���G���X��C}�"�n�g�O2 ���d���eDA1���5MO:�?�BC���vl�޸a�mj��N�@<��Ӗ��9�F��hL>�%��/c�f�K��H!l򤶵)�țd�7�\z��5uz�A8Y,�xr!����ُ���_����K����4�ΎϹ�"�8�*�v���%M�=�[ZF�;�Sc�G�z�J����L���B��^������H�K��/[�c�?�O��N�'/��5�SH=���5J�x�1z���{	�m'߶���aҌ�:��~�Ta�?g��}���oUf�d�ij>�I,��0o�����"뽥� 	#�Gw�Vz�WoB+��e�����F��$�4����'��D���2#��sH��I$�F;yD*�NS͕Jzt�p}��%�ʠ�,����x�g�ḱj���W����v�!\���3�N�NTDC�:���Ε�ˁ�f�ra��\'�H(���9�&�U��8�+�K�����"����`$yDG吹��
f��|��M�Q߱D���Xʈ��n���ڔ �	�(r��K�F%q�U�A�n�����!�HH��'��
�5鱃�*�����]Rp<����vВUп��OSx��Zh�0��p�|��s��7{�3��8Vڠ{�P>��d��40���qb���V�W��ŕ��6~��J��Bvdt~�v�G��M,-
�ָi~M���9JnR�y3t�#hf0�+�@�a1=7�1m�
Q][f�ǀ<��f���7�؎F���� P8WeI��?���cN �+��VsN�蘃��e]��+-S�m����fT9tp}A[�]G�~xP�j��̴_��x�&/�9�h$v5���F�8i��xM��_���p&���o��SW�S�'I��1<"��`�g�B�S[����jW�W�{FG������.������I�������\���<�e�\R@��x�׮<4
�4�_\D^\�"�����o���{�/O1�::9���t�<���(,�� ��k�˲�����%hDDDF�S�~g{�l�u�$��w�7,�Y4�KP�)���5k_GD!�l���{�N��G��I����'��G�ñ��p�8��b�Ёr��t��K����VA��G���r�Eh�����2���l�k/E�(���m9��L��q��������H¢@��苳mg�7
����"��A=��������pp�a�E���;;=5@h����r�����ѷ��z<JY3qmQ~��2��y!4!`I`�t�%�H=Ԙ���J|��L{���)Y�z$|�H2-&ڣg���{v
|�ť���M�L���/��C���u��٢�$��α��[� ���PE��P�w,'�;l�ZE�� �0�=��*e\R�C�~�5,������(O������B(c�񡶓/0rj��k��
�s�o����D#�������^u����@�I� *)��ЫU��(�U����ꑃۋG�kpk��Ж_��wH+/���D�T���Ͱ
�Ɂ��P���fK�	�<��PhV..�6���k��x��ejj'���k#;�t�5V�g=�-$h��1�U9��t�fQ�����Х�y�b/.I��+5�9�.��g�f��h⭃\I��\k׼��JT���T:Au8���i�V����	�h!�ZTs����g��r߄�iZ>�ڑ�[z� 9��iG��y�N��Ƥ9�{8��.��,���j���IB�y��)�z�0XͧgRQd��x��u #��gg���&|$SƏ8D�Fd5QxC�����J����ί���͌�c��1�faQ��׈"��ơ�`{�X*jo_*[��J��(�Й�q{��20H^��ˌz<�����u���㤃�������V�g%���Q���b�Q�X�}	�����ƶ����Z}w�X ՘	��Тhi �\��?��j�X]]]��j������w��%&�1��Y�ї'1/l� �T�@jm~�I {�����p�^�pDW��wU����: � ��_���� ����2�E�(�CV��0xob�J⥙a��-��D-�I?�6�A�"�>�e;�f3���"г�g�Z}Wu[h�hx!:�T6�:��P<�F��w���K�"�]�����Jg�p?l��J��r� �*+./�J\Lx�~�K��ȴoOS+A9�7��kJ��"�H��K�>`�>N[܅�͔��h�������e�>�^̘�C~%B���P6͏��ʰW�Nݞ�lm�w�����iii�|�ܓe�(v�	f��" �}��j]��읗�*
���~�P�b���;���/��v���~.`���9�H81w��z�?�=4�0��1F]��屵�i�<?@�9W3�{� $Z!��Q'T��e� �7���-T�� `��|w��ގ�

gl:��)E�l�+�ҳ��\�i�DЄ�K�b�;�Q����S�"p/zã���0R����6�l;!�G�p	n貂�ҥS����D+-�9���W�j��ߋRc0����	=`������^{��f��#�!M
w�I*df�x'���Wiu���$`lgW�i�D]�ca�R�t^o-���c����ޱxT��w�,�Ā(Kƃɂc�T屳`pۛ}쪫�3��Ǳ����Đ�[����7��0p��A��nIn����TX~^��K�;
`q���SQQq���Զ�RA�%�#wa�.N��"{�h��R�7]�1�:�թy�9 ��p����9T3G<&s�X�W	Q"-���Q �b~�Ԏ
�y�ݿ��G�KÏ:/�P�9J/^H�NR`G�����\666P� �/_��<�������8�C�i��`4_Y	C���aJ�㓒��Z2jgT�o����$����:<)��ff�/U�d���6?��j��;�>0ߚJ��i;�iߜ6v�e�ʻ#![�Fʤ��'��z,Ť8)���H� ~(��*������:�A�eSA`	�$�
��z�B�����a,�^l*G�M���|,� ����x�ډQQʉ)x�h�Z��/i&5�n>�\\��ʏF+Z� ���]�wX0��?d���{���Y����������\aa'櫊�aԼ�/�a� 2�F3:.�s �92rr�OJ����d``��k�1�L�]@e�dʨ��Z���4�|����/"CI��0�H�xNiN1�rx��uh�ճ�t�� ���N6<8f8殗wgg�d ��H���wIHH�fH�BƝ��Ǌa9`V�,`p�*RV���x̣�W-� �R7��j�f�Q=�D�>1B�m�I���.`I|֯h�����HJ0�KRqw�?���g�)��85�>	�f�����#i-�"�z���<�ڳڡ����?Ĝ�O,���+����6S�;���GƧӂ����ue�u耍�)�\I�	����H�d�l��O0,/C?���)MT� ��ʈY�I���C21��|��ț"3D�?T���xc�8�4�*�h�A��mr���-�8��3U�oj�7M��!#�>�`�;m�Q�-�M�+:��3jpS��� ��`��{N��~,dhJڣ����v!V�2��o�(��Vr�0�4j�Y9��&qO�)�X/�9fC�R�!�./�	--��F	��8�lD%0^b_�)���N'&B�$]���n;Z�^�fI"D`k�{��'��y���)��0L�4MRA����}�E	��ƏX%�W��}n�*�0=1��k�*}?ġ(*���r��M�k�������<"�{_e��Awa������-֏�� �|�2� ���TP�y����m�}�.�����p���Y���"��sf�[**���;��M��|S��H�q��~q?�GQ��|��:��o��RأRu��j`�G�f�D�5�r�R����˃����W�ڴ�w��oC�SU��0��&����tX-�rJ"�S�_8�������U<R��z�Xl_$�,.�6����|hϦ��l�O�N�x�/v8���si샛�Yk��9sdf5� ������JJ�o��m@�뎂/�^�J) !�/�WWgq��{�S&�w����A�-�=G��P�|��0]�9E�������f�a��?����HH����䫠�l�h9�W4�V�b�-�Hݷ��Ȑ5R� D�.�,E.\DKC�g%�B�'\�tta{q�,�	���(�쬬$�Bm�w$Ix���\!)�"�R{{��L���v?�=g��[�/����Z
��I}�%L�
��T��S}�ǧH��W�Yz�P1�j���N�k����T<!!yl����\K��mw�_ M���G���Ǵ�o��.6I����E
��G,�l�/JQ��b��db�1�֨����Ѯ$���_�b�V��������z*} ��羨�8���$i�&E%2h��t4����K�$��\4/_��D^� ��r�W��J�c�� /,J;�g���o�߈չ����Z	nȆ�7�$�	���/�
�-~�-��\MU-���'j􉕹��q�|���ݼ4W|���:��g����C��>1��0L��]���}e�Q����W_�10�F5T�6W��5vc�7�m�V��q�����AT�7[��W���(4����-�5�X�ZV<��Dy8��@w�\��u����H3�z���:�֢7Ԭy$���o����K��}��"��߬��k��j���s�*�Q��VN0�[��f7f��a�����o��[$e"�t��������1����Q�G�{�J�h*<�u��P��<E��f��)ð��A��Ƭ�Y+8�C������@4z@9i�E��:����9vp���[�@�5~ �P�';?X��/�k^����,�j��]��{��`�Q�1f�*Olu�FI��±�.\ZҏpրWsM�" �,$F��kx���!�z}��M���ᷨ0��������Z��mv����0�$
Ued	���yz��&�$�6a��C�''����z�'qiW�^�s��>s9������c�X"�ӏh���}�'��tA:]�Z9�,ia���+�"k�ւ��p`�t��b^��ׯːMo.ۣ[8��c�S��c�k�eIY->L���wI�d�h}GT�$G�I �hvq$`gg���s�T��7�6m����<��y���?R$,*�{�>g�G���[Y���9�F�����vçM^hJ���a޴���u��^kfTTA��J���co����t�H$-ҔB^\��؀F5�s� z��},�	Jr������K�����
ߧ���׷�3He:�gj�O���JT�����L"V��s8|2��r��l%�+�i�j5 Z��n�45���F��xzF���0������2A���\��jof�'��J_���Gr��ٛ3���1��ɳ�0��2:��wS̸�J��/^�+fQҵ��0�����g�C\1����0_���9A���F���8Z��^%��a\����yt��SL �}#t�������ۡ��a��E�5'���6+���Yn�FM�k1=7��2E��o�6:GiC��)���G�xؘ��>J����'�G���7��YF�Sȋ3F�Z����"�ֺ���l+p���5��,������]O[�EU�@�TЕT��s�ʗ-�A���i#ɡ��r����[Ak|�g{��O�f��D�a��V�p�(���o�-L�w*���ԾF�P�:>����!������Hi8 �5^�>����8�� 11Z^ê�jÚ�H��O'*<��[|��19�-\�����Q��������OB���d��}`��:�C�fi�c�����|�C��(�,m���p�6IvZd�mZ��.P���8n����SA��UCn���P����/u~���P��o�R-lEm������ `>�/�,h��͟����''!3��E:��4z���3��EKf
���c33�W��,�������C�ya�4�q���7���^s�d�;�Gv�}�"<�
+�?8��=��݋��r�XBf��t)�qv
��~t�M�:������(o��z�>�&چ��o�?C�g�x�>#ޛ� 4�x�P$�e[D�_?Z��yQ��T��j�á�wq*�m����G/�jjb�Wgf���2Ԋ}<Gh��j�։�4�Wje���s� �,�P��7%do��w[�}&U��$����c=��eƎa`z�w�"8��JMM-}q��9P�U����uuBl�X�Hܺֈ.X��(�*��߬�ǰf��QS��_��r��ޝ�R�P�P;{�b�
>�����_��)�Ą<�8Y\A ����� ��)�5��N�U�!W���m���M XAq�'���p3�����:���hV�6r��]nVͿ۸b������]'�^7.U���0�g�d��?�PI�6v��s����}x��rT�xbX7+?r�Ux���?!?ʋ'�<���Ϙ�<UBZ?c��ĳF$��~f�U�z�d;��[W�ƒޭ�{..{{�"�M*�F�@�U� }AU�0�dZW3����"6bjʟX(�{p����TB?[#Z��g�����Xܦ�N��P�˓(k�c�BM�?�X�ٳT}T����}n���0�B�檀�ʎJ��)��#t��	�?�Y�XYyq�zzdn��]ee��Nm4赟�۝���v�G��������)�e��C�&�ӧ��f�����+q%9~& ����݄��O|ݘA1/3�x�=��S�tMX�rG�kͦD�`AA��k����1r
&�-&"���տqr���;�̄����9�3k�#v�@
r��q�?�!T~��d�X8Z����Ϭ��5�\?�%;��f��[�B��{g�+0��̌�\���Uc# �E�]X��ך���t�^�/$�i��rE�'"&���	��m�EyC�s��=��ȥw��}<�{{|�������»�,
�*lz+'L}�3�}ܫ�n�V_j�Mݭ�_mˍͣ�V�?�������}��d�]P��O>>�:�~l��+��W��
g!շ���\�ѕ���'�6$���.�u���Pղ����ɹ�
!����>�i#�n��rFj�O� z�B��$S=*�䝞�L.�����ʑC4�=��d�7��FoN���q���"@�eXo�)M��}�g��P���u	���/����*��a@�K�ߜZ���Y���Q)��Co�V̖��#h����c�Ʌa�A�w��ͷ"K�nJۑ(!\��ߵ�o��)-��0�]����4l��4�:6��͹Y�ز}���20+���T�ԑ��٨�6��F����	N��T}�ۿg��$R��+�IC�~	D�r���!���s��R�|��~:��ۿȞ<H�O�9>k�(���1
�o`�wh(:��Y���'zm3��L����
��+P��45�o��=@7u��"rr�%\X����KKL�q�ag�~�Хm�O�������	��%�/e�|(��j�US#�W��{�j��Ko��>��J�q(��~��tqv-����}T�>��S�9�̟Ύ?Ņ�+�̲߳/v�*��Y�G6�����&`������I�R�EE�X��',�Cd�<�R��;J}��&/���C�Kk�F!%�uw��.��u�X���������5�o����Z�E����$��ih��9��cf2N��ַ7�p4f�#�f�+.>�F"�L��o.���Y7Lr,����kX��h�Jik]Hf"����6w���ؔ�!�t�����6x��0߿�%���n�5(yC宐�sM�D�A��^��,/�3����L��e�X��\�$���Z��	�H�b��3?�8���z\X�Ĩ<���O\R���f�|�oS�5�6�Rq_���0�g�p�=������sb\�H��1��U���h�/���	H�e�����O���\��P`�cՐ�t�&,�|1��e7YR�W,Ԭ����hz��w�_'\>�.��S�T�+b�F��_<�R؉z,�q�T��3�Z����B�=�O'o�f����?0�=e#8�R�IArxN1�.��M�+˿����S����e5\�+���v�UmI��TMǟ��bT�߱hK�=9D�L{�/}����=�.]\E�Lvr����o*��j𨿰5L���[e�M8PUXy,-��!�Z�]����p�a���%�F�e/o�Nb��H�4�����wm�Κ�ʿ�����L<�{Ȑv�`�*�V��鐙A_ '%%���딑�@4̾;Uw&ZY�G��D�R�۷���\13���RL\���)j�.\A?`}yЧ�+=9�]0�d����R�,�� �����%kTC[P+�R^��x�����I�ȿ:�(�����A�����p*'�MY|�O���y�Zi�i'�����YZ[��δx��,���A TCe�45U����$���xZ�=G^hk+�cV�&�yOz��̈́U�p�g�!vq2��O>.�dy��!1��l��8>&��m/�	�H�)׬�T���[����}�
�a�>Q���+�֘�!�|��ݠ+�}L�C�{q��{~Q��!�B�{Q{P�ͨ����M�I�}F+��JpϽ�s+{,��ˤ�E�'u��R����
�&�=Ir���U��z��Ώ��$�Y���֊e=q�@�;�^��7���e�����u�5Ej��R�].��s2( ����.�tO	D]]a/�654_YCwG�޸�/8\�.#*�8.�A\g��++����s�w�?�w�#���L2k��bZ��/=rePN�[E>[Fd����G�_<b$���C�}#��b~C�\:�D�{9x�֨�5{��W�E^��H4 �We8Y�n}�k��V�!=��>�QAmk�<��Է�HGէ����x��>�Q��RdX�v�M�-{������<_E��*�,d��>bJ��!�����P�p��z���d6�nzj=����	-����L[p�A���,�n��؂hY���wG�ւ��:y�}]��h*<U��~}i���lꇄF��J���Kpī�l��cʮR��^�7m�EE0M͡E~����܈�y)�LmbRL팦eh�؊�o�~�ׇ������xOs�.�_-hccsc�I������vh���kjg9�b��ꠁ�m��pk�Ny�<����5c'���S8P�32g����Q��55ݮ �%x���kN�n+Q�+��;�PI��';{K+���E���E5-������\2(q���B7p��eV-�Gh�kMΗ��/��PK��9�`&�נW��1)�xa�_��X,mrSƌ�î���F/*b�3�_�����I	��w9��c�l:_���(6�o,hlLs󆽙�k��u�}�QW7CKK+��]�����-���k�􁄛��'go��lW'�A�����Q��Q�p�k���r&�%Z\O�Źʬ0�xD+@�%:NN.�eM�����F��hFJ#�3�'��02�)��|�C�#��J,��_[$�i�9,�t�8���?Σ|�i��JQ�o����3lO��b*-Z�q.�u!���Z�j��8o�b}[6�x��qS�a3�2C�x�c�c����?��Z��*�T�#��������`G�'w�")�1ȉ����O�8�~���{��$��ep�ӟ�7�vb��|^�{Z:���ĺ�[�B٧���M	K�.5����l�B�8�����6H}+���:F�T
.QݤWXW�q��;yu~>�>'(ʰ��"���rp��j��oa���o���s���#R2��ѺA���z8i��x����Rmj�k0!"!9���(�D��TC;�A���i�fS��$d��\������H�F� .�ς]˪�{�0Z(_�����ߤ�(C��v7Ec���T�����X�t��Ӳ7�$~<T���-�<c��c]h��i���S�w�MU�6��̻~�F3�N4����d�܎��}�����E�<�S��B�~b'���W��.�lD�����A���dT�����(K	���������<q~�"0�s���Žjkgg�"+�S~k�(�]�Ho�����ZLˀ�Ȏ0����2��b�ޏ���v~��[w���?�ƆmM���]k���`��p\���MB�[����s'���U/�����B4[a�����e�7�2_	��@�q}�KͿs�������T�uv��~#(�5 4�̢g8A��(�4^���gh���� t�CV6}�y#��1��K�K_���|(U噯S��D��n?�f�RD %˩�q���Ax\���`7��;������\��k��������&0,GʦW���\�����Nwl����-t�`�6����Da�ra��a/s��gBBaS%�+m��\?�5��88������yq��2b҇lz=؍�*��@ɟ�,�O��j���-��;��QZAyo�)��Q�gX��{qBޥ��=�Z�L�$�t���r�u!k#jS6�bl%m.M-f�|����h�ѓ(�f�����K����H+jZd�]F�啈��4(�j�v�+����/�RF��*=P�s䊑p.���U�% �3��9��i�&�oK�y�Y0S�e�j�+ 1���tY*=��'5v?�y�^\f-�bQQQ�2+��L�c�)� :"��ć-����)9'K��Ժ�{�˾�L�O$����j-��żE%O�#���*t6�6��b�"sW<SY �͍#��?�~¢��%�\�������w�^���+�U0I��Br{���e�N��+��it�|�?-4��������}#��2�a��1��X�m��8C��&�3�è�������l���+���n�k��"8hS��Y���
@����'����>̓�eӃ�������H�b�סqS�_�=�J`U%:
.�[�.�0��>�`�I�����A�7�#b�	��z�+z6��U�����[����}0I� �'ڔd�������6ԥa
T�T���qQ��<��W����X�q��>�h=�j!���b�����m�:�w�Κ���T��pyzz���Yj������k�����(�z�g^��B����P�lL���*`��%�qa������^�j�[�%o�?��9���0�]q��F�h[X$��3J�k�?� J��ե:#�5e��¢"%������`��u'��-e5��}$��I-��[���Œ�>v�D��a�"�X�Q�U�����~�W�8tQHw]�l��c��o�(s�}�7��S-���"����mi��O_~��� �n����A��/�����x����33h�����P���=P���뙝+�����b[����Y�������U�ʯT�7s�c娛A�Wkv��T��� Dp8�_666f��!��&p�oMG�젦F&sK�$��f��Ԇ���8�}��)�Mh��3f�߈ű��*�+�>B�,�oy����y�����!$h�EQ6��X�Ǣ<���f���<�&MW3,�"��t�@Y�a���ji�]����Vx�i���ezG�L�LR<��̚%�#��oX�z��o���/��Ķi�J��?��f��;�	���G��G쫡��u�������t�;~�?W}U|����J���:���T�û��GG�hhi'��µ���"4]����b�J_G{6�E.,k�Y1��ǶaM^�K�ƪ��+���[�`��=�],��?Iv���&������L:���k���/?�U:�(�H�{--&m��`�-��������Y�u����ڟ��0�)��ŗO�V�m#QHw���&/n��WK��y،I��Z��f�P?=z�1v�@�eX��J�/d*��K�y��0�S�>�;������$�8m���g<�~wF)?��$&�ѱHO�2�0%�Έ�ܜ�&~�H�dQ���ڷQ��(���ְ��܆�ݙߠ�B�&�����s��%a�9����k;ͱU�?`���#�z+�	J�Q���İ=IsS�kO�C@�9�c]�F˻�x1X�ih�<�_c�$ck�h �{�����޾��D���Mٽ�W��W6U���0ք����X�3"���s�P	��>ɰ;��:��h?}7���ȳ���d��Une8�1>?���MI#�/)�6�.h�='S*��:����6j;;�Y�c���w��������!�~h^���`�(ौ�sJ V�fC	��UU���|�hw'�p��.D�-dƑ�g����^�Z���vpqeU?C�p��_0���lJ��{���%4��>�<��fZ@$T|�G$d8���r����h���4�qHf�lOL�ǜ2Θ
��۽��ܵNW��"BC��2�i"��5~}�?�q��N���F�B`�׸���ܜ�|c��_f��30�:6~WĎuϑ�'{bGHO� �%�������#4ʕ;U�E� �	֘��6���&���0�ϥ������&�x�b�Bvz�*+���K.�3Rl�7=R�S��׊���,l��ª9�/��s{x�b��DaPƳ�H��n�EVS5�A#�bۏ��^��]���44/`�/ox�5�l�l�/���KM|�=�</l)ª��K�xm�h2��0��Z?i(|q���rXM*i�f+)#��#�Y�L��������_k��#����J	w������
 7�T򄄄Sp�c����E�־�+�[�vv>��}'+{�i�(���w|m�y��!�uhC�0�r.%^���I,�,���Ϋu�ݷ+nڟ�RW'&B��G�GFF�t�M�jn���li�9�🐀�x�0���e�~�c�ޜ%'�ֈ((��30��C/�ť��J�˹W�_wqâ�|I��/	��Ѽ�v\�4�s�'�z�J.T�SF����Pk7�N��������B��z����/������)����Ʀ1����_"��?=e��[�������$�A���_�:���)�ܭqca�s����PrZMPY^u�}��ه�)�Ra��0���E��Ǩ�����Ӓ{54A��#�;����p`7��Y7�^�3J8kY��aܱ�Fd^0m�0������Q} b?���>#_X��s6���~�f��d�	l�Kg ~3G1�XO�;j��G*JQ�JT�UVTuJgzyO,k���Ԣ6���� ��fJ3y��7=#�� ���֥��y}}}�^Q�]U8��&4��x$�[\E�ˁL.��+ě�W�݅�uڮ[ݩ,y�2���f�w������M�`�,�<�:/� �Ӿ���7���	M|@2>P�}�xB�ß ����E��&����g�.vf�8B�7U)�4����K�p��H��\��$)�p�[o�]���G��`��k���C\��p��/�z�31�p�.�]Ύn~����c禋����#�����\Jd�MO(���x���.���c��4�2����:[�U9y���1���ivy�O� G��p�}/��O7�^]Mi`b�U �N�Jo��j�)���|��3N3f����]���9���Si�b �^�G��?s)�!��vy�N��� ��/�7�)�f�E�W|�(,!�T��Q���"$x-���� N�>����ͭ��	~���������g>��_�s�7"O�L��4�]
t� ւFrU�k���mf�I�َ};K���꩜3[��mK˛X:M�Jfb$�u^������bՔ=�k�ī��(0�y���B>En��E���Y�#y�nYBBb�QI^>���
>����Ӊ2�� ZU����Ae�p�7�3����Q�X:������O㴟C�G��p%��ɐ�-��ߊ��aQ:W�u���Ѩ���+� ���tQ���x�1	Ν�^.'�}��#�q�{�W�L�4[�%�#Wڟ��i���w|z�{�g��)&��i�����}aa!�flo�~��RWC<8���S^=���;�ʔ�.�%a�A�zVP�$:�t�#߁8\���!k��#��c���F���I߁~����b��"�xهFθ�����4�S�}�j.��b�a��u D��I�Q/4 �?ȰTkj����O(����m�n,�m2u�?
�0>����M̖�ݥ��F�O��٩�|�\[�/�Q7����bnΆ������dg6�&�$�Cn.��F�����(��q��jGwYBރmB�M���6I&�i]1X��۽l��6U���� ������3��bT�T֡�8��ռ��.�Ykk�	)�wM�qw�}���>�rH�=eK������TŲU���ȍ;����)2��g'�C����v���*����I����Rݭ�P�F�eǶ�:t.�Hw{�6J��^�����I��3���#�x���W�:���!��o=�{�N�\�M�9}�g)��,o'�*f/�����b���?[C��@��#����\����P��ׯ^̀� Ϳ	�*Q1��eS���xV>>F���eM�fǚ���z�r��q���5VCXû�7Ʒ�SS����] .���lK�,��$fpM>���b��z�uc�]�;�	��7.��xZ����L)g������*(�1߲ߒˍS=�x��P�!(G_[�b�X�haE��$8G�HLD4��?��+�-!%&�_W��d���ި�g�R�+u�r�=l��O�xV�؁�EW���2�$�i����"M����T���)^G6p�3���K+����A����X��ƚ~<i��RRbkX���)_~�@�gg���r����������Iq�`-J�2�kӻ��8LY\�A3�F�N��/?*bH�S���{:���<�V��d�����5��|\��]%���3F��C]L׹AQ�C������_���ONb�h��}x���D?(�MeƟ�L���>������y���x��?	X��ɨ3���1��Q���Q����;�J���		n��n���Tc����KWi���q?	>�����t6�\�P��T8(�Z[���!�:fa_�}6�'�_�0Nؾ�R߽X��� vʋ�3�o9���]E�Y���{|[�kn�* ^�Dc�g������Tjd:9�CDBd[��S�dQ��;-����F�F�J׌x�]�W�R�
-���sbP��犈Xt\A��0���?|5EGG'g<���S`�8G@L$b_��L����)�A��X�r������Ab1�hD��:���5:**O�ܺZ�W朩ͦ^�g�9c���g��c�_wI���i��4�}f�U�t� X=.c�	e:HZs��ÔcQ�7�S$x���+����M�'/��=:S��|9T�VE5૗?���9bi�B��S�����߆P�0IB��?�5�1'1�����p.K�D!��X�M�h�9�Twg�)A^,��풒�<%����I:��85sS ������0��zI��>�]�A �:��i����s��?��n������F̘�q�A��>~��?�_nz(�x��p�o��d�#�Z.ޫ�HpС�������eH���%�X�4�33Pm:��A�'F��8�j޾7��T�!o��y
��x������zs�*��Q_V���KwHw+�ҍ�4Hw�4�;���[D��D@���n�s��｟x���{����k����[�߮r.J���hs�r�S�>x�uom��%���ڢ�����I�b%ܔ"/wo���]��ݐ��@�����WgQ�� � 7�\,�\�_���y�r�ں�0|wg�#��O~�f=�D��0��T}i�����oԒ- �C�����]��A�z����~���}#񄞸P)/|�$�:6Ɓ26r��5F��f�(�Tv�~� M���#�r�����s���T{N�N	0]W=���j,��L��n�qۜ�e+���O����,**��N� U��i��q oh�$�,��i�2"��Ե�p�i9.���w����2�3��>F������9�o�V�8J�Ʌ���<���s��Z���b����+ѷ������7�M|Q�lE��,�|�27yt�u5X��8(H�ո<�zF ~�e���?:&�Q�8�z��ێ�?|x������<\I�C�Q�yy�I�X�$0f�|�����qžuPE�	O-S��%�ԇb�va9派�ATwww��u��o0XҨRr=Kl8T�����al��$�SڗK�2��$�=j=pa��
��� G����S#����C8D�+̽���)�?�i��;�Q�1�������o���7�,%�&���s�E�ymθ��l`pY60{˦�AV�M	 �m�ȅ���x�� ,��d�as��s,�����ɦx���T
�b�7zR�#S��vJ}�;����E�:����-1��ɯv���V=N�������~l�8���5�*�ب�S��&O���l����<�|��-���]�q��*؛��n���;t�8=ߍ_<~Z�>���ˎ�<��$$r���sY���������RO�p`N�|� n^t��xF.�(�pm-�(���[ZZ��soT���
�����^�mM�Ӫаl�U�E:[�B}��ӊ�I'��|+��No�\�m�4�z?�*̥TkW�E����e�x��n���|g�j���h�L4&�%���ґ�7���߸a�MG36�1��_ρ47�Kd�G̿�¿���i�d�h�^v��8��W�5&���I�����-7T���2%-ѵo-�f���K���'�8��&��ւ�����p��N�I���ۇ�gOn�,I�}����8ᓖlXt�5f�Y;+(�dn�I�M�VS3^M�66]o�i�}W���l���jcm�H��<|���}~^��Q.ŵ
�S!��{�t�	�] �o�ʗ���aeE��(�!0� --Z� �/;jgo719ɤQ{���̴����hB�/�Y�Ǒ��QK���6���eL���}+v��d��"��=ea��7���/�i�y���&;5,z#�4CƷ�M":�-d�\|�@L�dC�N)�^��h��Y��}�� ���f���D�����ϯ��+���Ei�ƥ�P��V����M��?��0�����6����-��5 �Nv�R����.�-UM���Y����q0��ُu���(�,��g���W2:~���k����c=�� u���L�<:-���X{0���y�JxN�9Mi�Q�#|R� ��|{}��2�R:�H..雍����}�8�ar��Z��+lI�98�BDL���r�@�b���Z G�%�}ʷ���f" ����"�3���m�/,/�2~�*��HJ�y��f%ءq�#�h����z� "�.��e�p7k
��'N�-�Y������6���L���y!:;c�Rlj7A��؄�SH�#�W��P�h��9��w�h��W��r:������ry�aݹՅ+�l'ä�S��E���M�&uE��;��Oh��WUS�R6��Am�%�9��H��/8?���>7����,q�^�b�_�jyI������$�P�,�0 T�.HcUl����W%��8Th�
GmW>����O���p'�"� ��zN���i��E����b~.
k�<�Si��|U�R��? G�\�7x�|�ˇ*��\8DIX#x^A	�[��
�T)1���p��h+���6��b���R8pPКp	0��J�����[]���M|D��h��+ r�u�2��:p�%��z��7�������5�h��k$B"�[���@�ҫ�G?'&>��~�?���	VL�}
�V ���J����F�ψˮ5���Dr��y���d�b�哓��Q�H�y���4�6�\�W�=o?��M������5jw"��]�,��ZV��b��D9�����_ p�sr����� ��F�K������n\%��[��Z��ӱ�{��g�!:�Z�����(r}]O{G�� 
xGdB��f�b��W���������%�;��	���fZh�ܵ�n���-�'���m�Ե*����嵍)	�@�n@�gGή~��6b��/<h-TI
��9���om�Pû3VS��S	���Mݥ�%��(1gK��&%��#��'�3d�
���}%��j��jF}��?�'x�+��ph�������Z����q����� T(@������D��qlR��.�4F:B�����IǇWn Q�[�{�d�wfn������*�lW���B�+�˼+��Ys��$�K��jŌ ���<#���N�7&�e{�)�7dwDa�u] �A%ؚ8)4}?0�*Q���(z���\U�fβ�ˉ����ي����O��~��/��M��`EEEC��'S����%˦���[[K�����&W�#"#e{�����|34
��_��S�w��w�#	�-|N-8m�Q4zy �z�wL��˓SS����.<��A��S��S�G\Nnv��]��EE;C?w���J��JÀ�]��c�v���nJ��W�Ot�LP"�bX^D}Pi�c���+�?�j#�]C�h�!Ý@MN�5sr|�/4���a
�KQ/�sy��T�������W��X�����8>ޚ�g�YN�{d�{�8�qiy	���^�` ՝�$37�L����?-D�|���pt4:N��Ú�Z��^��kX�v0W�'�_C��XpU�a�K9ρD^v��]_�������D^�;fB�X ��WN���j�Ws���$��9
l�%�<���.O����� ��~�I�7��gӒ�s��vh�Gk�;�FF�+�М1il��3S���<���jH�/��~u�������k��U 0S�h5F��E�6��*���1��yB���'AX�Gǋy���Q��s�J&�-^޶(&�,�7�i�Θ#�9�"���BC}���c2<�Ŵ�@�1���{��M��l$����ߤ&�^�<i>Q��J�� 4_W�Z-�9�&�M���<	��j
=�]iv���ʴF�g
�M$��o �,�Bc)�
Q˛dTr�W֯�-;U4��+�����wp��Bm�#B��b�G,�����"�����PĐ�_#yЉ���C��Qm�DA����&p�ji� �ێX�/ci���M�i"�C:�~[�p�w��y�~o���0��SS�f��arT� g��� O��[Po|�bX�֦�kқ~]¿@Z����G"�[ބ�P��6��nw��d�e)����ĕZ�����b�����A=Dӹ��m"9�m�8XLl�qQ�E�FF�V~`ع��l)e�5�RB$��5�J��q�"�A?�
,��e�B�͠yN/��J6:D� l���W{���R���%?�.i�!zc��l�U.�K̫/68/�(�&8Ω���p^�6E�VD�Ȟ�dD�^���E���N�_�k7V�e����@�-�f�!̯�=u��������o�p7S��j��/�����s1�������ZVV��6x��v[Ż�����F}}�E��䊊ba��+ǂD_�ʬ�}�WT�*�s888������Gs���Ns�xY��^��c}��a%��}�Ӂ�C#甁΋��8�絡���X\�
H�b�ă"��̩�#�q��{�Q����e�ՕT�wr�)-�b���V��F���p����B.h8})+�W�^�6�����'9�bC=�C<�च�a�yN���I�-�c�_k�W�"m2��c��$���S�����@Ͳ��A�-��]g�Y�����sԘǢ�A�>~����6���ӌT30���VZ��
@��q�2=A`�Z�'[zz�ܩ�ѻ�Mb��\z��
�k���#X�GŖ1j�3er����	�B�;{��@:��(�����o	ƌ������no�m�4��@V��>m� �
		�ͯ�a��������VAn�_:;:�4�#~�����@Z�JY�������5
,K�^�)`(0�*�l'c�����(V��^����~N�������4p0Q?�`���UD��F�buVv֞�	j[�q�� ���h�����~���7ng��o�5�KR���:��-�������f����3$���%����E���~K��fS��W����ʟf3+
�=����TJf�������L/E���tq��������~̈�[�%ԃ�gJ*����D$U�z�N����ٴ]��vJ�������ɨ��+Nb�������oM=��.7��1���˹�Gծ�g�V��$�R��!+Z�L��b�B>��h ��l7�Ja��<>Գm�ü'�ou<R)����Gk��?��������߱������On"������	��Q���2�r3QZ@��d�����#R!�31)����VE�S�!���ŧll�#�f�z��/��F������ a���A��7	��H�\����n(��_��Y�-��R��+��*�̡Y<kϫ%�H'�(�wG�m�`��gլ`�Q3�KFp?�Aď�5C�CP��퍑�a����V�&F ���G�A*ʜ%�@cT<����҃�^>1}�x���8���vh։`���_����Tvv�����h�M�Q��F/ү(h+ی�θ�9��P���iKQ�\"%l�j�_ )�@N�n؁��_T0�m���U8�V��r�2	��=
ք�K��z��v��I��M���h�]ɣ�~V�`KA�C��_�h�,4,s����U9���~���#�@.�H�V��_������frb"�H�M��i��{-�E������B�����A�d-M���`�Ϻ��?�X,�@M�cm�C�]����?�s˞jB�t���8M΃�� �[�oFA�T��Sq+~��݄r��eL��z���K��E��zG�=��ݖ�:{w]
TP\hh�fH|W;�2��A����ƍՑJ-l��&X����|&0�ڃ<���$�S%J��L/��̬�����Үs�D�S�T6$��塄���ڥ|bb	�����9�7m�#����i���%Nv�#�~fS*��rA�p��eA@��5yo�� r�V+b�l<�Z%+�6Si�l�/�{<�����%sk�h>�P:�Ғ��8i<�XC#.�O�=�Ɇ�ͱ�����{D�L���tB���۫��$�V�D���:�}�����p,�Ef^ �5/�i���œU�S��._��]���j�=^7Oa$��~
yWQ����t���L����-9�T۷u |�%������_qV��C��.�����I���A�٠��$g�a�=*^��%B�u�<���TZ�9Y�:�!��H�mu7iJO�8}��Q��e��v�FƢ��Ѩ�3!A勒��j��eJ����f>�8�@�N#�7}���m�
y�Y_q�"j=W��V ��R	�q���T323ihi��ˣLR8� o�He�,��]�5����d�ol�%�+�<�5yD�MUPf/���vj��o�w���V�/* :� X]W�#)*�<�!0sF^���n���Y�˫�Ha��С#Y/��_��E����n��a+s�cxR�ُ��3�X��/W��Z����6r��u��.��$���٭U���#<}��8�����	�}�JH-�v5g��h@xG�C��hX/`B]GEP�涳���!���;�	��^{ϕ����[��ڹ�pQ.��Rלl�͉3�d�#Å�Z�i��V�2S�/�!a>�%��<��mm�N�Z~;?oLZ�E�n�?��kūP���s��Tc�����{2����Ai�B�D~c�g�.�a��� �ɫPBf��f�d̌��θ�҃I�v921%��_;�]#)H����Gl���_Ƭ�J��G�{Þ5�k�HP����u�3�P8�wÞ���
�Դ����q�E��ZtQ��{g���|��,ЦSm�o��D &��2��$�Z�P�W�r��e��]X�s�%��z6`�
g�E��5�=/��̶� �׎��Cw$��.�h`�0m�ޅ:1�mՉ� ���� �?���;�G��z$�ߗXN�2��GV��X���2���s
�^+��%�x�b�=cT���BD�������'����\���[YYY5�0�l�K�rpo�Qq�絷l��b|�F�G�Z��"�O,,Pk��n�k���`���S���vw}��n�*���L�ؗ�j_�f���5��S\�l�xD�َM��?F�ac��Z�����:�G}��r�;�do��Ƿ����ǯK���)�-u�Ռ�g8zA�z� �)��P�֟ȑ"�ޜ`FJ�Kxx`:�e3���@�J O�,we���%l�5����s.�,�7<>���u������Y�2~��$�|�箘����YԺ.@��qǟ�P��������R#ka��@��
9k��#۔{
�|R�������g��Ο&�5�����[��#�6���լ��[N�[J��EyX�"K2��!x<�`Oc��,8�a�-ID� A���dA�1�K���w��5}u��/EŅ@He o�������`���4&V��Y"�:�Dߜ�2`@�L��?ܜd`BW��l����mJ��D�=X�`� V	��yW�?�^CS,=^��7�K읮{���.�����pVV�݋��q�F������m����^�x�ۓQT�a5�+���oM��M�&ۿ��8wTT����}�� �:U9��6�N�N2�@2Iff���7��S:u��-��x�7�]�`;� M��ō�ZEUhUG��+o����屝�\��:<_ �7���lDr*�s�j��0S!�t$}g�06B����pFF�H�Y@�s�	����D��iKK��ӇS�|)�R������$�5P���̓^d�8�Y����0h�pX�E/
�����ο>��3@�\��kj��׿�������R�$�c�����k�� v��E��^���n���˘�����̓���e�L��34�[wwMy�ԾrL�@{q'1�'[l��Ƿ�x��K�C&%]D��Ç������}F�#w�.B��So/ͤBK���U�o��\
��)Ks���!�f�g�����}W�B�lq��s*���֜ĵ]���2b��d�6R��K�l�ؒ*M ����'�x!����6�0.�J�]c��s�6�O��gr*�Jh�H�R��3����Q�=$�̊Z
p�r��px���%��h;��
�5s�!�ܬ�T�C?{�3��G�$#��j�R(�]]��?�$�f(���![��>`!O�tH���h���6��5�%�]ĸ���H� gW���%�ݏ&��,;�v? ������E@Hp���	�	9�T�����|w�7S�-����P��7Цɷ���*y.j���SSSQD��6����gy՘nʦc$�4^.�M��k%f��Ȧv��Z�C$�K� ެu���q-�U�w
�|U�/���)��	���Vu����;�ߡ�l�?Z�C$Z�:��{���&��<����ĐC#t=��_�@�E�dH���EX+FDF+$@�m�r�8I
e��@y����h;[��0�?;ޖ2hE;y���������H��c�!S������"&�9�x*2/�|�D�z��C���a\,Vo�����ܿ��+Ϗ�w�a�g����k�4�I�W��= ��[�ȥ�&����a|��R��p)�RK>�B��d��\���f�3{�FvN��$��A�%6ۿ��t��H���]��@�q/�|�(���� u!���X�c��L1����w��q8hC�||qwz[����u��eA��*��;��uU��f�wܩ*�<0��ϯ.~�锠b��6��y�FO���b�c��Z���e��Ҹ
�i�]*.;��Rn�P��V���\ D���#�lY�$�}ؕp'Z���"pS̐��Tn�R�CP�{���qa|�3��/����VFs�!0���PkiCz�0m&�$L���e`��F���Z���{�Z̙�x ���!����}�k?Ұ��O2�vg��~�4��5S��RR�&�Pu���R-����!���_|��z�&gC�
q�V�����:�%�$�B�N�!�߿������y�FI��snO[Kݹc+D��#O�4}@#66
$�!hV�bƲ�b�����3Ȧ��H'��>ѥw|G�N����Іg��vAZ���ܲ�:>!!�� ��c�AG��H�+UiN�V��9m{�hO ���3nۙW�w�Y�j����7+�_ۿ�k-������A-�� ��P-e�ITqؖ����d�
�Z0Ji+�JeSNh�~`D�����m���K��xx �����1���,Ǥ��I,͜�fTܙw$�<��D��,ҕ�⽌�dȮ5eK	Q�iV��� W���
�Y��jnG{�����?
}s"����A.ٔ�'E5�a�O��G^7f������ɜCU�F3|[
��
������� ���ta,~�-����9���Ѝ�)�}A���n�z=?���(��]�MB�ܿ�'o�]w��N�D�^^�+��[���C��Dַ2��J%���L��q*:MĂLii$�B �Q�E,�)��f4����'�O]6�a�7�C�� .�y�x?�Y���
H0\�-Z#3��8��4�e]����|&m�`z����F�W�"����8��h�	$6��?߉�J4�0�� b$8�n%?�͙�j�G"�3emv2D����ȾD�rCAA�@���W96�3��OR�����=r&Q�{��Y�>�|�|���"G�k4��������
y����W�M$Y��]����=A�t�~�nhn'�@�.��]t;~8Yjœ��/z��B����w�J����_P��O��P��U�JY�Г��4��4��O�bO�n�����S ����U����	�H$�!ܹ(W�CܹL4u=}�G~Z�#��=%�O�]e}���jhQ�)-*A>�����}_8����na�B����#�U?$	[��՛�"��U���R�$x��آ &�wM�ߎ(�����@R0�J��&�������)�X�6wT���o�*���c7����L���-<	e����!��`�Йʶ���|�1�QP��*�w<��w��n�<��"�aw�77�D��Fv/�j�^;�կł����*M�)�	*4��.Ov�W y_�H����lk>t<�	[�}�.�h��w�ݳt����Ǧ��&$�uƗJaG��i���_Ք�.�5�.k! �����ߋ�M�3�q`X9�z��mE2S"DT��`��An@^:@27��W���4u{���O�^������g>���9,@��%���.�*�M���^�O�9T�M���ﯷM�FMc��JMu榃9u�*{��)�~���a~J÷s�����dڣK,�S�c�h�@��W��ڷ�&������Oz ڙ���?���4�Z�uY	���
��P ]Tδ͜�g�M�S�_�����䗓��	�xp5��/����nH]_-q3^>���̿^	��{tE�Gu��OD�����hM��Agݩ��<����K����g��Rb��~�*�aO��;^��~)[gg�p��\�������W�[�9���Յ`a�3&u�$Q"x�$�/o��"�br�P��;P���Z��t'Ƚn_�mG��܁���H�	�p���$����O[E�@C�s���kf�_
B�e��-���������32�^�9�e�J��6��U/e��)�g��fm����jy#M�{}���7��>.`������l��������2-d�e������ϕ��j.Y�l�=LK�y�b���	Ż�V4���LU&D29'���mX�i���8�T=5Λ���0�b��Cn���L�X��7<�?��k��ÜZ���������8����kC��.����i�d�,�me�ap)�yƩ��?@��@��d�D�#�Y�1�G���Έ\�:��6���i]�l�7O>Q�O��H�s�h�G�a\���p'P}ާ�n���F��$��1]Ȍ�`F�2�U�[H�Y�n�h�.\���p��Z�qߟ�����/:No"r���p[sFK#�$�[Zg�If�Le�\Kk4��83���S�g'��d��$� #.�$����~j,���}��,Q~'�A�^�ߋ�T|��*�z�s�R�t�<�8����V'�/����_��B��������LoМ{�%&8�����|�QGUlx����6�B�VY��I4�����
�9��yA���JLl�w�/k�'wP��u��HK�K9bz{CbL���ʯ01 �5(W���Þ��8]oe��P(�O�?��T����s�ڽDiR��g������ϻhkonj��8�N�D��p�%���1R$�[}@�V�zn^�4o���K6�&����U��V$k&��DDm#|���Aeg��G����M?��]4\�a����=��<q!7N��4��P>?7�i�)��$�v9� ]e�W�8C%��COV�]�*���H����{�V��k-�L��_����·P8貘ꭈ��"�̃��٠�ƚ�x��.!+//��DJ��;�`A��OD佞G��ng�G����0пTVT�r�b``� ,K�wO�ZnQ��Tyr��*L6c�;�r.o:!�[x�9/{Q���o����W|�;���''�P珝���1ɕ+ϮR����<$�~&i�:���|���o?h�=)��h�����T֠��H���,l؆k�]h!e�[�����8��χ�+��e���M�Ƃ�7�/��Gp,�x��p�֑�郶�?����ӄ,�z���3�M1��2s�6I�WZJ"�s��s|S�Ü�#�{�m+K[��>7��/�.�S��-,��v\~_z��F��J ߥ��q���q�=&���1cc�l�;+��AŖ��e�o�!�&wu������FH�ڱ�<��w�ݜo�a'�B�?���>�t��n������o���N,�tm	���o-�����9�Wq���,%i�6�����Ϸ�	�G\��H���([�^�����]M,�����Y�� ��#_��DRo��jXRs��#Ņ4��7	L^t[VR��j��$�{2iH�O�$��ɽ��4���:X�#��,�aԼ��>�`�4�~��>�g�;1�.����6���	5�ɼc��X��α�H�o����8M�_f��.�4�L|�n���MO֧L f�!�j�d-5O�������ӽ%�~��'�mr��٬Ю��ʖ�{�͝NYY������";��X@��[җ=�bl��Ҩ����y\������y�W�x��2�%7W�SSS���{]��F��60B�?���-���ګ\W<h&��k���b��B9w�wmq�?ℙ˔!�Kv�-%�����>��k���%���C��Y-�4�{������������3�d���>��kHG>���Y�}�8��tP6}[��o�,�Կ5�؞��t�I��K�?���'��Ո�����B�t6=E��?��n��统{R7��r.��L���.U��zu?x�����M�5wvR�ǦUh+?/����?�a8�77��\ݦ	X��I�XD��[��;�_=�z�	y�4i�\��;4t��W% �W�w�S��}p����9>f�����ũrt�����ۑ7Wr��eѿ�����ɞ�9�]W�7�II�Lc�0� oo>%ҏ%�;�p�>��+��)DO~��.������ma���9�,�\�K�i/�\'e�8��G���1�f�������p=���~�����15n��� i-n�F��X��(u� ��-m2rH���z(;���M>�M�4ퟷi��ttt�4�ϙ�Lv���*k�����w�w��	̨	����R~
T(�X�<�w<�(���L�������m|zr|pRVX"-�;��
P��kH`G��h�^�m�ER���E@������C7�����\��?4DQF�>70��Y��?�4�P��_��o>��zr+\��kZ�/���-}��Hc�wAT+�}[���|�g���c�#���ix�B��v�". po-q���Rz��3�h!� ����ŕ�%:�]�)|�;Q@��61�tr��#�"�V)�dH�{�3-�Ѓ���跷m|M�	�~�u�*C�~dիc�Q	J���*��]C��"��4��M��o�����yx�\�S6��/�^@l������p��<r����5rC �9�����}�I^���R�Z�t�xd�|o'�<j^+��?���`���i�
!%N�]	������m�}�=�$b����L�����cL��*��,9�a�[�#-?���\��$���-��������4^''R�	=5�X-0X^F^��͈�f+���Ɲ��~&��HQ�/j���Z縊�����TŊt�s}�j:���M	��d_f���<?��؈o�Q�K1�.ΒN��8�~ ����e�����z8�6F�L�cZ#!�Y���@L���g���(rd�;IY�{��`�j�
�� a�#C��黺�P"��=/s�]H�x�}M'�][y[��Rc����ze7��[������z��������B'ۮ� �I�A��|��q�}|C/xi�@�Lw}R�"ͿN�K���o��� �$�>!S)گ��Z{Y��S�   ���g!��+�v�3�j��XiG��������}�&�	��%g!�.���@�q�9v�;v�r�YSJ2��'~}��n_�R�/�j�����Ԗ�p��|>�Q�t��=��ǘ�|Y�z��М����g�{�j^�Ɂ$���Ǐ.��'�G��c:�������K�n��͚���8�(_N,�����϶a�-n��_"����}�׽�nV��ҭ6Ĕdkz~���:�7T7�{sIu��賛��,���p��f����v��м�&��&XXxU�Vdbw^�W�ᴴ�4֍֎_΅��7�|d��1���/cA��B`o,����/�zeL-e�����BMxo�"u�؊?����wv~��҂ӄ^��[���-�=��Bi�1g���2�/=;��kk����s~ݕ���QA��s���%<��3t\��-!�W��>*r�V]��گ�=��B��o1CBąM,��,*&2��R�����2j�H��]��B�Z9�kD�$o#�-.����ȧWAI,��f#��c��K�o�xm���-'�hoDZc�o9�&0k]�tv��E���u���� �Bq��q�L��8�L,�[ȧ}��J���l�;��L�	zT�w�RбWc*�d��O�{Ĩ�����λ|hj]��PƷ�kx��(��Ki�ߌQe�v���j�ꀔ07���u�*B��4�4C����!���(Pa�"���Ob�O
�}cP�yx�Z�!�g��ը�u��kB/�k��BJK�ȨN�%����JL��[|Y��'#����u���\��a����V�|�E��ө����Q �QP���sMZ�@��D\0�i\�z�]Kv��y n�.L��J8W�M�^���_�4V�����#L{J�:����ߊ^�C�a]��ı��𲓕S�A��O��p��q7Ȃ�:��;<�m��C�����w!-���Y7�L���ӡ�O+�t�.ƍmo0>�o'�f@�[rM��w��yw�o�m���_i���O��_J*T�E�R��'x����Okm���\��˿�Ͻ��~*uU�v�#:%���m$b���nv|�I���'Շ����hM_�U���P�_�2�f�W��8k�����p����O�2������p��cu�}>�ez���B����l�aӯ�4�R4����zG_7,��X���%��i�ϗ�!��h�"a�>��÷%�L�V��E:E��,�l�����;i%�m���l��H���V����
�Fj�����
v��K��3���CB��'�#���t��c���FG�$���'��x�`X],��!P7�{�J��Ґ�M7t�l:r�M�n�o�ܡ��+,ߥ�o���=1��� �l�D��4#�. �ފ�e�$��-QÛ���1���vY�Y��߆ sM���x�U�>������Dt���CN5jQ�rTG-��}z��@K��AI�z�Ź2A��\kQ �C�f��P*��A"��u��0�Vۣ���(+�q�c�zY��;N����5\#�X�1}�*-�;\�u5�z�C��H`I	�ٖQ%2�����գ�Rb�Vl��+��`�1j�W:k
�X1�}�v{~�v�0�]��}S7}l��P�<�E���1I�{0Z���r,k���W�\�T�RR��/�U`i�����0�0�vD��]���hA��!V,��u`�,�w�����[�b+�6��JK)2h����	�6�ۢ�lw��.w��>���d�?EsP����ŵ�c�Ku)�����U�i�cY����vE�h8�0�l��@���#�!�Vk�$Cu����$wX��t<`�m���D0rC�X�y�=7t�����v��X�N瑲_o�!�~��������m�
�Q��ӦuQq��c݉CY��ϓ��AI.r?�i��o���#*��.��]��2 �x�@m�x�X��#Z�-���z����妦�u�����!����]:И�w�(�颥o�R �XP�S;��t�ȥ#�.����ո �'fA~���4���G�u�t�"�Mw��<��[�;�vX�t��_Br�s�q�
����_iɘ��8�~�ۯg�;�)���!��Tno4��'��#�W��7' �fmp8CI��M����
�5�3����68��n��%�k�m��>��u0\���g����0)��I��{[#�lb&&��*��j��ػ���Yb���+%y!e��#O�&��1�mU�'������i0���,No��9L�.��8���p2O��r	%��H��@<AEt�l��>�>� ��Uj�uoTX���3;--�-ѩr��i��l��ݟ]�B�����Y�|3���d�1�'D����"�:9��y��F������2��lȅ�G7���}M���TF�(�tp�q�.�8og��׆����S�'�K%�4�_0�c9�ۖ.�-J���ju��§��C���zϪ��1!i����W=+)ET'ݩ�>�G���ـ�/���ue8t{���91u���g�ETh�{P� �89R6D�J	F1 ��H^��*u\;��AT��Bq�����"�K���ݺ֟�q-�����E��/2#����L���O�H�<?֖��G
[��`���fϴ-���-��v�A��,�ɖđ��nc���qeW��3Z�.&Z~��o$`įxٳIy%�M����]I���#�fp ?ic���S�o�2�n1�Z(Vw ��������K�W�Ϗ�{Sz�X�Y���G�m��3d$U����<Dr6:;�tJAy4�S.�t{\�ˁ�{D��`�)ؿ<������9#�py�������Y�h�nM�˛;f������1�����m�&�=�8�UNY�:v�G1 s���R���J���n�c�l�͊����m�^�x�9G����n���6��>_���6It3�O'�v�rn�6�V��a�vى �C�����J��t�cu{��
2���~n�c���j	KUK�M�k�=�����"Ȱ���H	בm�������q**�z!R�T`$s�qm���5o��Ay# 
�$p��)7̜�g��L�p9��ٌ����䕋I����m"�lZ�a_�C���׶7K&�H�{����M�;����Z�k=||�״�5���|B����]����[����Ƃ��JZ.�����	��X!�,r�2l�I���
�������5�z��N;�Zi~��~<j�^?��n8�dɗ
)�/#yD�xeA���9���,��rs܏�Q���g��fj.B,��;/Z��ח��'[�G;yANr�Y>�V��&eչ�3�x<��̫��!����Uru����5�a3��r�2��>�S^��I�i�$5�%��F_�X�ZD�\^W@�U�d��q�M[�]��>q��4]��Qo�$C�oB�O���o�M�v��4y��]��x���,'-�u3s󭉠��=�H�e×V����pH�έ����@���)ߑT�,P�t�C��u�`6i�.�f#�e�
��Hy�拰F	��ޏ� 6�-m�t���(�KZ;��~�u���B�5�`%8A���	�s�g��E���ѿdDx���o[y���c�޽J"���"�[��5+/
�IƲ7�s�%W�T���'"n��ӊ�`�)}e"��L|��C�$��ݯڹ��.1���`��V�x5N�yÿ��^I䢹�h�ʨ6 ���+.%��{q(����RZ��[�"���݊kp�@p���?y$ٝݙ�I�X߇+no/�%�x阦(�? �@X�cpN�0O��Q�ɍ���(1�{"IQ�1�f<���Ҙ\�Q7�~�.�}dP�Ӷ������ ��U�ȟ~������n�IjP�URʱg[�	��֡)�S���-M��*'��|	s�#�*�[�J��5wt�Krn�5����9��lj��j�4�̅b�pލ�$?��[�p�>�k�M�5�((7m����Zq���ѵ������d�*�_�v�ѡ��5����r_�Y� �Hf�f/o���+��g��bUunɧ*��a�1$�b�l=w^Mӏ�@�r��e��jUqZ�8��M�O�E3����ڌk[�L%��d�d�&���^vlD����Hr z1��M���e����mtI��1�?�(l���z�
Z^��f�p� �G��qݼ���c����4�$R�n�0�@e�� ��~��a���P�M��b��{=����z�0�0!?<�R�a7� �?2�{��8��T�ѵښ�����*�[	3X������U�@�ʷgk���=���7���O�k��D�rs��=���T��Ӭ� *g��2ġ���y�	x#n�.~s��}�Lov��Ν*��P�q5~pq�tʹ]^�0����B���E�~�M��5T^�4$��x�rWR���@�A� �Ռ�]sa	Ju�_���2��c��*9IeW7����iX:-����3�s���	i���A4��Z�-��f��ץ���A�e��ݥ$U�°sy���| �O8���5O�zt�}���uq���9�G�6�b?c�°|��n�r(���}@��C�(~��]}U����, ihˠ�-3e�h��W;CX��wrS'�?0��d5�e���1��i�U�*�艓�;���BH�Y� �`���KD�T�Dղ��+�
ْ6�rB˝RC�&x��h� ^�հ���|	��1#��-���~���{��H ʡ��U&�VY�*��V�摾1�����C��h�ԁ�@���f>���[�;#�y�)P��p-C\�:p�M�!�����/@ D� W����hFt�spV�!k!q$��~4Ҙ���ӓ���O��U��^:v��j2�Y[���3U�!9�g�:��s�p���
Ȉ�V4E��>�?K��$���tЉ?a2v�K%K�W(g^RbJU��'=Ω���$Q;�C0y1�rn;���]��U�qa�>�<���~�?ME`����'�^!KV%/yu��Bj{'��Zn�+�T��k�z�H[2e�AM�b�9��{&��;|ee�k@z�n�4<�
���W�O0~�������r��#w�_j�s=���t��8~<M?A�0�E���d���ˤ�MMl�o�B��*o�.^%u��`j�k�Xњ�W�A�u%�.���(�P2\9�_gO���y}#�$�\iGj
��#��b�l�$���U���^L���Ok��&�'��q|9f7ne�����6in��F0V�*�*�{� ����TK��$����5����>�l9J�4 2�=~��	�xA�Q�[*�;s��k����ڇ�x��M3#W�3\�O���/��p���+'��I,,��	�pູ�e=�|z���$w(�඼�FJ݅��̙'��VO����� ��g*@'2�R>��.���5l�P�E����\ѳ%��BE����B>ڻ�7��Y*�8�����-��K��R�X�nk���ݭH�8�1��A��>�|��+8��{���u?�[Q�0aXЊi�:���6�����;�Zk�w�����KRJ�L_�et�7qIڸ۞�D���	;�hz��:�9���V�c����!�$��F�~/D� �B����3P�5T��+��y��!|W@��};�n�z�-'#����W��H�ά˾(���q����G���HaD�_핪̘����w�6���׍�<�u_�/�y`f �=pC��R���wUy��['���R?��H�$��
H@�9�3�3��\4��ުG�'�f�<?����#�R5���,�e߯ºay��j��&V6��q����q~?w�\����؉r��P����*�¯GXe�Y²��hA��P=l��3F�_�=?� 	%�j�%04����h������V�� ؐ[-��������Z����r&�*���HOLA��7����ښ�D���E��D�&�(���FM��/*�F�e
�����^�0Q���,9�A��g��A�|V�}��\��5��ҽȀ,��'Ns�4���5U�|�5���ǩ��I�	�v� �~�=^����P��#"�h�e�����Z����w�E��Bj���m/SA�0>l~���o w�����[�I�}Z��M�
��F:��9U�A}%ʮ+3&bi� <�[o7��)���ү���z�T����N/!��ޭN��5=�Re���\z��?��Ϛ�%1�H�,�[y[���k�F� ��� Z�JA����Fm���O�Q������C�&s��w[�c�H�:��VƓ���6I����#�3�EO�!�Dη��TS
��M���X�č��m5���~���@�{]78�d���Y\�㖏N���H�г#�:��-��~�	:���[��-��Ɯ��53XLc��ɐ?}m2�Wh)7+i7��Y\���\5�2I�V}Q���l{QS%���UJا��k^
�7P�z53��.�ݰ�@�l�.˖��|��w�[l|o��CQ�������RCW��Y���^��§�zղ���qV���}9b�ɺ�z��2�b�?�"QV��|�x���?sJlg��3���*��:���ƹO	�S�?�IZ����$R��w�,C���0�E>Rb��A{ǹ�B�q���[����@E��M�ڿ���/zPn�n����'K��K�	I��0�� �����4��{,ن�z�#P]Р;��́��\��G�c5N~R��1E�}����@���=%tX䱵00/.��,TR��ک�<��, 2�mW�<�ì�PL1�h&�@C�Ơ��e��д��zXڥ�>�H� 4��I?��n���ןۙ�:ZoI9�B:�F��7�b�Rj�2������F0j6����߮�����=Y������'QR�URͭ��W}��~�v���}m#�c߷+��k+��#[9���wL��كHd���t��n��x����kP�1/�yz������{��I{�$c��<��V����ͳ�=����Z9a}�h�4I�/X� ��q`�h�<�"�^=À����U���@﨎�;��9齃g3��Kiqe�	��4\	I���Ɇ�e���"�%
�K�W���JX��b&���X��i�&���0]+����F�8��j�T��D�\���t3�������ʂ%���tku�.�U%��F�⤖L5~�"�{�j�m�u���v�E�8l��h�ޙ�K�EH��Q��k�Z)��
ݗ9�`g�~�0�i��J#Ң9k�
�����IߩÛ���MY�$N���%�,V�>�A<��n_g�����d�_{
h�S�X��3������8G(��߄�u�BG�*����g�����?�3b�~�\+H�k�1Q�&�~ �Nx2�Z�j����Ux�>l����~A�x��Li9eB��b��pe(t��m+H��-,�pze�y �*���u�Y�8�l��Z@_a���a4y�s��P?z�my�P�3Ç�LI�̎�$>�z�ˋ�2�P�{���$4�g�{_�d"�M�E��3ST�c��s����ڇ�mz\���d��w�u�f�)�m�KO#f������bL��S�P�]a;ć8�AB;X�$��9�x�z"��@C!�l�c��)f+T6�י��#��Y챯�M�_��ʫ˓pIn�W)4Y�3������;����4+V7T�9G�Z_u�1��?!��B�0s���'�r%m<�L�1+���C�w��X]�u� �)�T���]�	��χ8RZ���(�����2��V��������X[��,жh*�����GȞ @��@ڇ1MUH23ӳ�邙�L*�{�C�����	jVFR�Ʊ�6)\�*a�,�C���g����Y�.7�h�a8z�up����_�<�����&[$�ћ��@�A�y��2����P�������f`V��VG�)��H�ӯPt2 �6�%k`�x��a��������"���P�� �1a�"�0p�QQ�2*�?*&��u�6�w��F�-+=��M�g�/:!!NWp(�u6L ��w�������\�7`���Kاph��P"9Ԑ�]>QB�����t:��?�T�n�}�ϽKe`����/���#��%O00�J/��n֜H�7.�J4$"s��[�j��(�&������wWo��i�d_SmŘK(>��x	��{9�p�]�]wk�qpm�v�~l��h�~�=ӊ�7Yz������n��SЦ�~�_�:~VFF�����a_n
�&�֦ԗፇ:�F���0�U���0}P�=�.�����.��2.:.�8�c�����[g-כ}����;2�Zc��_5�q|���~�@Կ��x_5R_ ��$i~�-:��иG$�������T��[`���5611���ldt>3�s��f̽��`�8�`]$���O����K���G
wҐr��8��8��Z�z,J�Z;�S�	@�Ĉ}:��H��s�δ#�*��iz��ҋR��\�\�7�I�hDF�g���⪅?�e�u�� ��pN=���s[%%laI�I����������<m�3�q�]�:N�>h�y��c)�Z�˱011X;���z��Oz�z�^K٦AgDl5�w���p����  ػ��C�>�jzMv������~��;$����z�qE�|�[i[1��}z�r�-(�7It����t�� ���^��E/*	�=��{_�-OxӒ��0/���V�q�n��H���Bչq�nt�m�۳hz۹w7�k�j�M�.�Yþ��r4��$Tˏv�L�_���N���'�*�a��O�v��~Ń��}���0+<�V7��q)3!G[
�2%am��Š[|4&�OzI����?
"�r;1���ld}����i
�����L�*6�"/0â�����tŕ]m�q{��SMaܺ��}�)p��+3l��ֶ<���+�~�R)V�;o�-F{)_`�V�!`�5��PR�Ʉ�;�WB���DC=WüHx�#�j�x��{�C�8 ��M
�#\�^��"���W��w���'�AM��}�J���Nv��ѮWeb���#"F$S���ڥh�J~3I8��1`���'d��|�!Z��z�=Xyͧ���Ny����,8\�M@	������?��6ljg��𱩑fy6����N:�>��B|�'��T�Qn]�?Y�P�58	 ��^����`>��YZYa�ad�{�0��0��?8y;P�Q��&����@>���Q0�v3(���Y�g�}������n�p�M冗UqMh3���qzU t?`�&1=����s������wVZt�!�w��!!�dF8��Q;�.�Y��l5�aɣ�*`Ѳ�9J����j���o���w�O�X�!��O�T%	�7uw��]�U6B�LY�g�3O=��O9�,긗�G��n�U����,��a<�O|;=�[��&�f�6�V�'d�r�XQT�X���$��h����kM�Q�=��DVq=��	���B�p��5y�jnfzk�bh�hvs8�]�">GN0Cׁzת�M޷@�hr�[��H�d�:����ݒ�&C�Gj�-6�!�ٱR}�H�C���w�a�Tj �rQ�|�����%�Մ(!<�h"U�+��O�I��ǡг���n�=,���ȹ�mdE��݀���r�PnDVu��]͊ ]��I�%��d�ܘǷ7v@���u�gl)Ŝ>���M�q(S��̮D%/\�n�����A\G�^��u�HwPc.�K�im���o�P+� �h�'�6�9+�ʴ�	�n�SB9�@o������)�P�\q{���a��� 5�+�Q���Ɠ]d��y�����hn��[�H��3R_^揇�K����6�>
���f���d�����2�[�8=��NhD�cv:�����%x)̭�<'`Dh4�S>XyCeA�8O#`�M���S���
4�/y��xj��U��Ⱦ$#�?��'o6�� AS��1�� ��a|�5h6Q�` �%w��tv�l�Ql�M�Po�� ���`�|�(����V�~���X�Tyi��9���6^$�ٖ2#�\��c���S}�T>I���ܵ�L���t��p��
�뀬��98!�+��2 �^�`�J��TS���z�:�/Wv;����
�R�����	3�u4�`t2�I���ƣEZf�c����JWmtG��ݖ�l����
��u�� ��ͣ�XY�=�~_ku4�̓@���X�]������6�X@���
�M
M���ū`���^9)��D]a���W�����$��A�Y�_�!څ$�WH,��F7'��a��;9�ȝ��J�%4dV ��� ����2A��wQИ�.m�!�ݵ--�����@��"��fz��±��}�v}� �X���Ⱥ���!݈e��Du.�-��0�K�p'��5�9�W�>�o汥��(��~:�sB0l���	���,ש�m_�B��9v�Q,���w�~2�^�	�~��J/^��גώar!��PJ}r�����Q�.M��[��pYO�fbg���M�\�gPmY�(�58@��v|���xL�λ$=�:�+�qω/O�� �޳k5UC|�Z�ŧ�i�Y&¢I��̧l���tV1Ld}����(���[��=i�!��מL�rwr
��w��\e��rٔݪl�^���"Ë3c��ԚԷ�M���	7��Y��>^�^��F�H��q�lU�lx�f��=D�
���1��l���\��?1�n�dӗ?d,��OٳCB���\/*k�V0:X��׍������
3��-L���G���Ŧ����WO&k��qF������/F�xAA��eS�Î��� �9I�KX�F�E����̭�И���RWɪUqٮ��<G%8����'�g�}�	�`}�%���ݕvYm����&�ّy6��'�vSD�6��_�6�e%܇4,��gw�˜�i��߾:T�ť��lL%�/�h�kò�BE��?�G�س���알���qao՜�՜�Sg(��Wz��pLX�����o%6ި%��Df�؆:L�]��wY]�Op񌾂��?��L�FRd�|LX9J����ou��_7���,;N�Z�e=�˝�����9�YЋe2�X���a)�.cQP�8�����0X�&���ZJ�o�$#�;��q�'��z�N�����e�$�1��i���ַ�V?�oc��L���ZP����.^��5%Q�A����.�	���~�5�"[�M���j�X��JS�F|R���S?.���8;���	3:E�t���>�g�;�629�ό��g���`�����`r��*�����a�j�f�D��Q��&�>o��d�z� @Ru���à�*c}Z"ZL �/m'�7k��/��;�d�/��o�U�z?�m��p�ē�������෥��cҹo���P������=ղ���UҸ&U�V�3��첹=�r5�	�x|��p/�~S�;y'#2�Z�婯����))n-������bӀ���䱗`8k�I���9 ��L�\4r�fy#�|����0,�D���+����ކ�@�S{vqߗ���L\u({�e=�����ƺ��,0��#�ڑ4a��b�ҽ�'�,�?Q�-��y~�ѳ�fy3�X��]���њ��ա�	%��(3V�9�'�j�H�������ӪAd6KS4�.��6���)n w����vW�\�J��v�L�w��zb�[���=��5��\����Z;��A�� �P�az�ŹUY��K�����ԑ����(�#th7cαЊ9����C��;-���! R������q���Y��n��W�	󰷠�F���E�
��ɑ����?��>�oWEU69
"��v�U�_�z9&�y,�a�3������o�j]���ɽ掬嵸����u'���O^�len�s\�,f�>������P��QOC��\v�����j�)���2�K\H;�
���zl�\��^�a�Z�ϰ�}Y�Iz"w�KQ8�ְg���9'�R��=�$I�6�1���4�p�h�_���M��SʾX��A/-.jظ�����m��A翵�밇����߿�kR6��+Yf�mi��2�u�\m�>?����K��v��@�f/�zg$U�΁U��H�7k~�P����D����V�~_[�i�yY7J�����g��V!S�;&�Ɍ��Rx�B �v�M3;?X�"i/��(��ꤟ�8Q�F���P���q�Rx�B�*�ok��IDͨ�	�I�-�v�$E�CU��m��������r��k�۽,�s)tSq^���I���������X�[߇&�Q.r��LE������	�B+i;�'�"?�~Zh�l�$�7hiX��s���i�cŜV�WK\m���j	.fŉ��ڴ��G�������r/II�s��o_�������>;�UYҰK��i�=��
�#���r�v���KmԿi�"���?��ڜo��w8��(��$�w�o�X�����_����?�j�?l�d��M�W�eBd
2�����|���F0V8� S��RPc��	�:�%�P�h����v��)��g
w-$�1�#���g�!�ß�`��Ub�����ʃ~�?�I���F�B�%;���oTГ6�[Ҋ}z1��ADct�I�zb��d/���x�?�gg<���s0�L�<����f�~�M(~ڑt���X��/���ɐw4ɍ����s�3p�#1 �|$i�,�fb�p����r�����X(�7����o�Rk��(;��G F9V�!��*©�Gߢ�uŜ����FI�Ww�1֌��sd՞�!��jE�3݁Ƭ�=�i���M�7;����,�+�`�n,Y@B�X�t\�P>D�-9���eD�z��>4��G^������}�w��4�J��5L՘h�{�UŤ�.v�)����_���gaN�%{�s�|h�k��玤�	��*6��4��kP�l]��V[�f��Chh7�Q�F�\kF�t����6�߻�0���d�c������Q�dCgo1�0���垢?i�"~K�5D�֮}Drr���cL���ʥd�Һct0O`�@W���j#|W�F᪌���C���R*a
�۟ވ��EP)�ur�N����y�%��dd���Ŭ��ĥ�����i'V�l�ҁ�̫�g\�z�KC�T8T�1�[��4��g�T��Mf���.r*w�
�a�7E�ԃ0'�]8�&�U�;4r�=�n`��m�Z%�I"d,j��S���z�K\/�4��-���/����D���Vs�O#)YO��k��HE))1���90Ź��E]{}�����S���|z0F���7��o
�@���(��7�����}m��vJ���"��*o��<:Ӻ�� ����-@WU����i���m�n�d�e'a����{�t0+|���M�C�+����,�OQZ�|J�|Jد�:���D{Y--�K�� Z�:J�u������8A��A g�E@���YЯʄ�����
�uNl�*� %�(�)�T��d�Ǥ�Z\���1P�W_�k�R��`U�Ilɧ�L�M����||�wwR��%��߀�-����b��%�v���k�v�qZKe�O~.xm��� �%?�%��r^����`ܮu�7�!25C�M}�֚ �zS���3���n'9�`�+�.�O �A�A� xWr#�L���N%Iem7�qݮB�I��"�NN��}�^��?��NjdI9"�'���L���14?L���'t��\���D��n	I�3f����Ń���*G�܎�=?�C�zZ�^��ڹk�n�!:K���2�a�EWq�����0=r9~�l�b�!:�,��GѰ̹�1�t�u�˕}��R9�?w^4�����WEq��z�[�B\��B~q������R1"�ƽ��悩���2�����8��2$����.6�~0�O�!�|���g�B��˕�䋵w�xH�9���<�%��40av�p����x�!��**�|��R|L#�X3p?׈Op���Sa�%�?�����y�f��d��
H�_�#[�L0tM�;"%����+�x�~|R1�5�\5mN9XZ��t#�V^,;|��*{8��H���!��r����
���SԔ�0Jrȸu��:�4�z����p4�Q״y�v'�j�詉&(�5D+y<��Tܵ�(��-\��n���SS�0�B&U�__*�*�o~g����]�H���;DG�g2����� �S�N�f�0 6.��"H�>��gA;�_�6��lw��Z� �<�y�b\��l}V?�Ww4XK[��q�9x��}xZ��
)1���u~dS�������:�EY������1����������xd1*�u2] u��Ŀށ�D#�-oL�nH0�eQ�%/V�D��R$Xe��EU���.ƚO���tz����mY���F8"�}�dY���h/�9���%�Ad_4=��_��������j�f��l�S����ǧEX�9oG���k�CNLy��t٫>���m�)�2��0\Ad��NnI�q&4�v�	Dә��u��;,}^�`����4mB��o
��b���T�O��W��[~��N:8o�Sr
���@5,q�(�-���׊����G���!PH������J�{�Z��[>��+�^d��x�Ƚ"���l�&�L9�aڶ�B1������)%9֯�?�5+l������L�����Q}e�f�mk�}f��A���O���@�짪��t��3X'���Y�-%-iaI����'o2��ɚ	�"����gY�G1�:�*��\�/R�Ȃ�d��zH� ��'#���&�
��n����QO��o�Y��oܸ����p�񺉒��ٰA����Uo���o�������K_r�������Ƣ{)�)յ엕�D����x��PZM5¹���A���{]U琛�.k��Y��[L�EJ�J"���1��������cY#o�o�Z�>ڻ�$x���PYhͧd� mWS�y�]a�l*}��4K��~��|�����mp���1�͡+@]�9�xI��K}x���ѝ^���������?a�3���<���~_�S�g`��Hĵ��Ǔ����X�w�9&��@�\p2�ڭ�a3"��t���a"�����
����wVк���#��py������km���#��k�Z {�_U�a�����|8bA)��cxS����Y������
�Ο��~T��J!��Z{�3���u�]3*Ѭ~%Ir:����Q�Q��LÚ�O43;Q��t+����޿��S����GN�m����}��늂n�rz%b����-X�̣�C�VL#��{b��6j�"��kh�@��;+�E_�77ۣ!AT]Qeix"Y�}gJ3���(ꅟ_�� ]��8�T�4���>�(�{����! �X�GA��O��򼒾��{�Y���6T~���7|C�j��߶�����v"b|��?�L����~�#o4xn~1��1Џv��]~#�V7>��]�⛑o�S�E&�} wL)�� �����?��/?�u�n�Qʸ�zζϾp	f`Ĉ1{ ��G-|�]Ub;;!L1�;���>A�IJkn���[#��qm��h�~��<C&@�a�YL��㯑"h�"�U�y=�-1<�Ѹؔ��q��WF��<��鮲u�5��s,*~d�M#b������W����\�������G�s�"�Ώ,��]Qb��a������V��6n��e�eQ9��Ж'� ��/�(+��`�Cq�je��U�l�sd�{^�
���6���:e�$�����e��C���_�����Y��\/4��}�.7�[I,ʚa^%�O�'���xHER�rGn�;�o��q��ꅜv4/��>��30�������	�:�P]ln*�6{�M��*��ԅ3*���) O"��}*>ڹ��s z���<�PT?�O;t�7�$��K	!�t�G�kkj����O�Ao��ZZAӧҖ姨�����0��Y�{w��+�#�����]�]���D�wY�1<���*³PM�B(��0zA~�܍QZ���F���ұf�w�iL�8�٣� i�'\U��O��������lξ��~Z�3�%�o��;&��8�ŀW���2�
��������>���:�w���׃��
��ۦ6hPC�3+~�O��tN*i+�.����>�:O7h�pN�/-�0�fV8��_���Ѳr 3�����y�Y0�m�_�ӌU�������s7�n\eC3;�Q �GN8�I��V���݀�*_����,7=��0C��ӭG��r�NX��b�䂧I�� i\25hi
��.`�f�)�M�`���W�o�O�S�a��/Չ8���SE���t��<��]��Q�ɓ�����5=�!��5�d
Y��<��� \�$~���6�^�!�����f�FTJ�H�>�������C�ۖ�,�/�Mm�Vߪ��_).�J�^��T @���w�wa�v���V�iU4��p4�r^$=��\A��W�?<��n�(�����L���<<�b]���\�N�]/|U�W����:� 3-�)j�$�7����¥R��O���8u�t��W�D���S�x3��g<���`�B'{���i���o��I�!���!t:, 1���+:'{�B��P5Anǣ�_=��y�o+l���%Q?&	w=y���H}�S�D��B��~~B�$��n���A6����a4����K���>ƶ}!�i�]}�~�/�|��0��y,��U�YO�U�}��>`L`p�o��a���2����8DAs���8YD��%��2]x���B�:����[���4��*�~?T�J���9����r�y��a�ʛ�ES̄E�P�d�Wʠ#���a_��З���%��ݬ��'*F�O��V�ft�/��N��_�`~����y����Y@��B�1_=�����3���=���䤎�F��S0�`f�5�5�K�/_�(8�
�"~K=R�zA,�>�e��x��u݆J��U��DB�l�T��7]�'�>�h78��:X\;cQ4Z�͖��U�,�N4�55�����ߝ�d���s�-���A�[�9+i�c�,��v��0�!l�v��C�i����A�e��o]��Z�RW��3���>��gʉFd��a��6P�̕�z.K}ǆw�P��56���_�L�K���9�^:����v�/�0���؋��~-�T�?IY�7-]���Ջ#��d��}5����̬ 4@����m�d��s�RH
� �m�l�y��q�NLCB-���\x����]�-���;���͐��Ս��ǎ�ac�\�̟���d�PJ�7���	"B5c?�R���?GP������aef��l����n͕�N��@�D*
��*D��o�xѠ�ס/�/�s�X��O�b�!���ء��̫��X��X~�;J5}͌���#��23LrW,N4���p��7E�'z	�S/Ad;�K���l�n�V��f�L��}8|�hU�i$��yN"�o�㻶y�Q*hkR2����%�k�i�r'��+`x��רF�$��gs�5�&d������7���<�7��Fw��<��
g���H"���rZc>ce�V�^��Z����ze������d�SW퇿O�o'����A��:�K��JEC�����鼚��/���}T���CQ��
yN�ǊA���D׳&�2���sEXY�Dq�,�դ-.�*֏�a�MD�1�+u״�����־}��v�9�0�F���{$��0e-�p��T�;I.���6Q���!�q��++^%D@�<�i�[�����v�8���B{,(���WQ)T�fl�;9}*����T�}m�h���A��-�U�YY!j��a�ZdS�;~n�r忭v�0�6t�^��\/����@��a���q�b��m�OwR�k*�ST��{����c����HG�V�wY2�s!����%!�x��ǅ��"�fMx��^�	�.�Fv����G�`/�Z|����Bٌ�����Q�h����2��Vg�{�0!0�0�u!2�Ū��}ꥌӞ�1@�3�L���l�R�(%Ďd��N���5cAR~���f�0#�$��$d
�V�1+^(�F1�����O��M׍V�9��*��
�(�,�܏��el�ღD3�Nۆ�Q���l��F��K�Ğ=�v����n�~�t:��{��8i�lbq1w&���	_}������<��5d.�����r��o��~Y�5f�#��Ķs_�xC�x\�d�&��Q�WU]����ä^��=�����K�A��sٚe?A����C�4>�����Djн�6q���GG��pa�?U��k\&s�����L�����mq�����6�hB]th��\:ֱ��7[��x���"heb�w��߃� ��!{e��R�Ij<>Z��Ld2��kq�/�	��esFq=�:)zf\R��p� �������z>Ar[I�m{jl�j���|���H��䜙{F�C2�j~���u��lj����fL�b����旤Ë���&=���B�f���K�k���=jԱ�v��!-^���i� O�_x?ɾ��Ə(�?0�1�^M�,� ���/V?�7"+!�@���p3��q�,~؅b�'AU�����PB�@`�����|�\�}�h��[8%���`�Ⱥ�����[��o��+tJ�=9�TY)�S~�s3�5X��a�o89�ǫJ�H�cJ�"_���3쳦�X[ģk�Ѷc�ic�=�(�R��1�R>'�sJ&ޑcˏ]k�=���� �=�!}�vVC�\� Ԙ۳\�� ���������q	Jr�+���Y/!�~v�ݐ��Jn�NA��w�6���#n��3��z�{`��KR��G"��@ìh�jq��-���C%�VVr)�XɪB�1\���O�h}ns��\��/!|	,�L'NH�G=��8�(�,����U#_6�i�� q��e�҆���1���Q�{�0z��7}AH/=�L���j��J�c}d�Ũ_��n}�s�U��w�YF����Z^�9�O������\�����m�i7��R��1v���_I�~,������&��yF�2�Кr����tf����P�Mߐ�4\�� 9-�ug'��c���*^��vz@�~J��W�9�����]֢�#�k.���Wr����Y՝��ǅ��2)]5��f8����q�J���i�f&�Z�/�Q��d�F��h�0%��d�}���ˍhKT�˓���d���x�����n��kl�x	'y9�a�EN&������?��J�Saə�E��ϑ�/�J�ZJ���Kp�m�:�Q���Xm��#�����瀷�	\�Hi
�'f=�on��H>�6r�5jNV{�t���:ql��[�#��^@�[�S���T��o�0��>e��H�IRL_���:1C��)����ź?����Ha:�o�@ĖB8�=koi����#j��.�%��ͰV�J��g`#ƀ����T�@o���%����I��n�c��:ru�dm�~�Ջrb�%��P�.A]���t�%�EY!F��+*� ��N��>`�0���9y�]�i���28-}=���Dz�,�b�UQ�@��T�8���0R���BERa3�ӕ�Ж[f�∀����T��i!WD���g��ddG��;)��V0K�.���[�Cސ�cϺ�	���I��?��0M-��D��ya:7���
��_m��BOX�6���ly���r.1�3&����ov�=5��U���#���f:q�~yN掘*[6=}���7�tO���X�gBKV�Ys�_����f�2m�,c{\7�٢�
(�xWC��ǲ_>#�z�<F�N\OA2=���|�����~�_�ٯʩ	u�i�;X�E���_���3�����W���K����+��w�x�EOe�X@�P��:��F�+��*�,,'Ϋ�sY|��57q���b~K�wT��I)��@2�z���"���qy�w#�~h�`�4H��[Ƈ#hl>����&T�݌����iK�����+8r)$��e}�ݝg���n�I� B�Ү����a����ֹ|�UG�Ɵ70z�l��x��͓�UV>�sLɸ۬i�%sF����^�R���o��kI�.:';�M+�'���`Bw���Qr=�b�+?/��M]y�.��F�%@��{%�8�������B��ұk��_�NFۍ�#�]b����܁A nc�3��f���a���M��a׫��j�.;��@���wwww�����ww�F�����;���y��y�^����ۧN�{���a�|��Џ/�]�����C�p5����H���v��ڟ�bD����p��_����5�ψ�Y����a��;TR �7�r�:N�yB8�����ڲ$��U.���^zp)r�	#蹯�/����O�af�O���
a�UZ��%�;W���>�N�]��g��!v��W��xk�b{>�p\�kQ3q�B1��~�p�v�{���NW
���s��~9slȩ��ϯ)��=~8�؀���O�d}�R�����o���DT�q���$|�:>Kb" {��(���p���I��\��k��iy���#�/�Ž�$!I�V�����̬OR�������Y1���ܸx��Y���m��X	�&3w gc�.21��xs٧3q\h��k���v;����Yo}������1@�E�T�'z�r����8J�|��>�k%�
��o><9����[��B��g}�x9��>�W��k2��Ͽ�P~�y���]��0a�`_<��C
���pg�=�܌,���_��T�~�(��V�u���$���<��@�ኣ6���?�8h��~@�1�p_9Ļ�������D�x/:�Yn�*��A��Q��@��ȏ�Z�x9�N31���)vZ��W%e�u�X��G6$�0�r���5К��u�vVK<��6�2O���_x�lK0��� �+⡫F��^V��ݴl�0ք���1`�����x��&Gg�Ct�d_9�p^��C���oX�D��(���3wcv�ұ�i*�-GV Rb[��K'̃�Խ�J�h�k/���tRe��7ܡ��4@2�����3.��x�Dβ�Y�B,`���#V�]ˤ:���PS�wH<�SM,�[E�7L��o}Hp�rf|;FQqhxr\�>�ٰQ����=��s������\I��`���?NP��X=���_L��u0��M���%�����Қ��q|$�9�9��8ݓ���ƥ[S��^'`��Ц���Ƚ� �=�ҫ�wi��no��2�d#쎚|�څa��a{�}7.�3�DS ��\L�|$��s��6
	�٤�=Cc��k���CF� �gp{�^�,c�Ѻ�>��)���C� 9P�_�n��>�$�}@O�!sn����̎���@�
f���4.�ҕ.?�܌��24��Y��K��e����z�����c� e�c"�9rRW��q��%�e���j�;"��~a8�h�r�N�����ڦ~��ό��II�G�{O�T�,��b��=����=mD҇��9\��EѤo����5ES���������.+�	�^7�}����O�����U�Z{0߹�_&�Ys���s	X�����v�K�t�RJw~TҀn.��@�y ݕ0q;U9A�NM�^8젦���Ѽn���ܿ�ٴ!Ŵ��W�3����k#�`���O��:RI�6�"���d}�ܞ���e��"��9<��9q>w6#����_1�^_6��u���ꢙlӞ������q�I:2o�o�|y�i�g�O��w}9 gv�9#_����ft��5��a�ߞ]�F3��u�vܐ��Wu^d�s�����\�5��^�従�U��9is-Ͻҧ� ~��7b�G$k����m�(���G��oK�?�{�4A�H�dI��֫��ނ��S=��0����Vu��퇇�-E��`���-xl��9��M@.`�U8I��|�h��-�׌�����R����~Z�Mv��gN���� �dHOX�)q(+��{u��Һ�0����g��a�-mKo�r��zDL�m7*{�)t�U����s%��@T�c��	�W�t?����l��~��.�O����}�	��j�4ɞ;l��H����pk���d�Z:�$��F��@� ��}_���O/|E�~^�i�\'�UK����o/_�}*������3'��>�@���P�(.k��}�
	�e���{����:�$m��?��~�xx�NX��@�2ش���C��A��P����O���	<1��������~�ъ��W���wefrxF^�_�<´
��MnUߓ7��rhk.o�Ӡ=��3��Y[k�I��2��ue�L�]�(((|o��H)�V}<oЙسP�c��x����/V�
}��]�s�ܡ���d9��2������b,����TH��J��4�6������V�������6h> 1�R��ᛅ��tAW�� ^�	�N+�ڑ�Y[��n��u�tP�Z�0�\�Χ�8�E^m/UR^�"Ҙn2�Cő�'�S�|��-ż�І�T<d��O(�'���r����?���=KF�/w�t1J)mZ�9��¨3�j7U�36�s��a��:Fi4SgbGOK¨*��[�s�X{���۝L<��)�RjncH���ۿ�+C��O�Ŋ�Z9��e�:�%)�͜u��+�{��U�Q�Å��|"����w;��z��d~�>�����	tb�OV�w"?`�C�Ң�-p�ihDU��o6����"8��G�i5&�kO��|}T�r^gN�~�2�1	(n2+[(��رD{�66`s���9��xi��/�
��fº6�A�Ya�U���ժ�=����٩$�cT럸�Q�	s�n�?�z���D��y�_̜*+�W���P�>�/C��X� j���=���+(��8�M��o���*Kai?Q/�h���t˴δvQ3u�ɂK� �D��DE�(�9wN����#��P����S��r~�\Ե��7K�xw� $h/�KnΣY	t��
�u�k��N䆍�w����֗:c9t�N��=���.��m�FA�����j3�Q9�1w��zI��,R�d#mO�F���n*�<|n�����6��p5`�C��g���a�#y�/Z�Qs�,h�-5mL�K~Z��w�����Fz�WC���6���o̅���$�"ˬk}/���~-���w4��ֳ���:�I��4��c�|[P"0��mUT��u�
�-�g W ��=w�i� m���*d,�pl��~U�ܸ���2����gd��x�,kJ�~-s�4���Hً�ǂϹfng���ݖ;��/F]�!�!"׬�PGf��.�dQ�I$�����P��Z},�?Fh����ݰ�i�Ț_��kY��d��H�������zlM���ZYڏ�4.����4@����l��
<�o�`�MC�PB��[�w_,,��s����=�M~�<�Y�ܕ}l�Vt�]�pQV�Ú2aS��,v"��з ��?�C%�䕀��1�moM�6��Ih
R��FM"b������N��v[��[uy ��`�##�K.�`����hH��He�̊�Ԉw�,};�	�tD\#] �h#2ڗ,/a���N��h�ۀ�]��h��ՙ"�rup�TW��`�!���6"v��"{�uv�[��D����C�'����N�}Y��z�N(D�G⦟��2WF��-���H�+�L�B�
�N4v6:�Y��*�WDbF#�q��>�O���ylk`ˊ���3��m �+�y����]�ͼ�w۔�v�����u�����;�!u��Ta��46��R�kk�W���V����z\��J�E���Z��燈�|��E�4�$�f�	��V&�7��Q����lt��_@w��K����X�$��R�J�m��{����rľ��O,F�Ŭ���NM\��h=U(tZ�!�ք��G9^��T�1V�e��ͅ.�Y\��jk+��Hh���Z@��8ZR6�g��ՙW���f�1#n�Na�`���ZF+��6`�����GP/��~���:��Ux���޴F@LG&��2$����m���V��Rl�^њ2�ZJNu����L7|�>��c�LYÛ}�������HZ<�V,�Qg�Ky3�P�e,jvys��UOO��`��'&��#z�S�5S�<�� D�y� ���]6������G�����~�.��\���E؅){��U+����X� �Fg��_·8��[��M����O��7�W:��F��I�i�Ǻukr�L
?/��Fz7�qȻ��I�`��z���_�b����u�3#��J�0a�V\5m`T�(��xnp\9ί���E����d���9\g�^�lt��ew���5!�=��t̂����� {�kE��3�<��>�79��	�
���F �<�0��{��:����z���+y���RM��U[-������������C�{I�%^��ܾ]��~}u��Q��	��i�Tc�@1�i��!�W�H��j�}5�2���dӺ,�K��_�
ur������b�>L�~�t��u�l�%Z_�Q[�e,_��hA�^��g�<�v3C�r��-_���(��Թ��@Hf�^FX�Z��a��u�8:�M�V��*��ؿʳ>�ѭѶE�-�/a�E{G�=0�����@5�4�[�k����*3����//x�߯�Ϗq$(�g�z��s�V��	0�{l��)o���K����!^u�j`�'��i 4�wB�Ɋ��G�KTM�~��[�Wӏ\oK0��i/ti��e���[�?-��9w�$��������.+מ i��h���kM�"+,�(���w�euF��՗��_m�n����̡%���k��cOW�}%t��k��Z�~ӘE��'s�����?3L��H�\� ��i\h_��м&�#�U���H?o#��(рmtT���/f?�U���!�ĊR�b�#�Wl+@�n���c���<��ͥ�����O.��wN5E���Վǿ��_���I�[�Ӳ��-�������_=��m���Y�	�X��l��?�坑���Z䆽2|�{8�����;�Aק��	�&?��%���|�t&<"��5�l/=��㤆N���a����}��9�,/%�����G�~1���\����3��aa��AU�|{�Z|��#N���	];h��R"���h"}VxX���V����]��[�5�Ԍ�r-|ߑ�AWC~Y��Nd�����֞��+v�"�(dń�'F�gN!�j��	�z�u`�jk7	��t�ƌ�s63S;�� �m�ݚ�qx��JM�~�R���6�<ݽՏ�0��a���fX�'�H�-m�>�i�I��G��><�	G�.�����z`-�!M�k���"�idW6����כ�g��.Y�[���vM"d�*��kci�7�/0�o������J��F����|���1k\0��J�O%VÏZ�р�Qcc�e��b�O�<X�#���d\��F��⶘-Q��!G��j�	>���M1��_<�H7��5��ۙ.����������֩�n9��u�m���s��2�;פ�e�D�J\t�{*�]h2��&���EM�S�ǔ�{&[������o^�E��0�b��v�]�x�j3M%#g�}����[]i��Z�}?I�7�Uڠ�>K<�֌��
E{*�55�*Z�����V�#]yjN�zzM�� ����u�����T٣2wH5�.Ǚ��?U�E�P�jCn��RPW6�#4��stk���s�z�/C��W�ݴZ��uG��w�~s~��*0��<��W�^hKl;p����a�Z���E��lʨ�=�9��n[1:�|$��N�'3�&�>.j�g�k5~C����I�}i��z}���.gYD�lr�δ�Ȧp׾Mc��IB�����Z�N�GDM$�����t��)��89%�M�:A��L'�ӛ$f>����5V����P 
����7p�^y��ח�a��9����ŝt�����	J�˴>`�"4�uL��j�@��j=��l:���,�_�h��3��k|��6��}U12�|�	����4%A�s�^��'H��K
�6����+U��)UM��j�:E��-I�q��+U��7�n3/�J�̈́p�]zJ��#&��t�b�12}"���P�׀�244��
�1��+��8� ���Ʋ-��+Pݏ����Ml��XD�b���H��d:/L������U��s�f���!�W�"��5}���=�,����4t�R��m�<�la9H���g�⢽������SP;1?g""ʉ��������EN���9�_]d���gs�JX�1c���V�@t�iZ�Bc�e��gB�UO�x�믧� 6�M�:���n��	�S�?�9Wį��'����N���O��.Zb�q���"c1�2A�Kp��*n�C](�r�Y�׏�=��,�;�w�?��& ���@�W�@�3��Su��Ҕ�y��S�.�V�R�S�#*uF��&4���ؚVa�������$�.kճ!H�ChϷ�qc��*��n�e�]�=�N�Y�lҧSYفe��
ֽ�xDm��
1!�PCő���׳$=>;/~#��\�/�~LwY��S>�!W{\.@s�(&I����&�^ՕAsڑυ���6|��˦���S�r�ړMkKNU��c�f�_k&���<��q��g^�{�%�?�u�����rt���R�������k�
�h^��tK���������J�Q�_���Y��H��^*��_�R�!C���_ސ�PO��=�A��NVj�a
��x���4��&(��L,�&~wJ!$�\�s�i�>;X�E_ߟ��?j��A�|�%�d��r&a�'H⋳Q�%���b��i#�Cv%Q�h��,6�k:�K:��y,}7}��k��Q��7�r5׶�4��]����zZ���2�CB�3������^��l�۱����AR������i�H��PF�y�-��G����Hzk~L��g�V��b�c���p��A"3%�`<(�1o5�ͯt�Kq��^�F�0O�`?�>S�����HyR���X�X鰜�_~^ڻŶ~(@ˮ�Z��HY�Vzk�QO�p�b.;���J�'�j��O-u�VMJY�6�l6m�"[�E��������׷���u�[�_ITs:�SK�Zv׭g��)�NYțεW��
�3�2M��P"��l��"�5|}�_��ea��e���~a�֬������f�%�� &Xm����c�=P隈���.4����?�k�
��:�`o&�v2=,Sz:q7U�Y�f�0�Ke��I�������q��z�Z���I��5G�3	5�	�鐒�9��x�#8 �>9H�=9�a��G0�Vmns;!ِ���ÿje��Q`�)~m2x�NB��ޭ�K�SD��jWld���Xbk��=DL
����H�#ͮX۹�$��V�I�f�����&�r�5�D<���ʭ2�h�^���Q��
�`����Ϗ����ǒ_p�48J5�최�b�R��G(-��Y ����?W(�yn���r�8F���[M[*��;E����
}�]"�"dC[�\Tݮ��+ϲ�>؞bV�^��A۳6ԧ/M�kLj�R�������Z�*�4� �8����1/���b5�J��(	�������_G��go���$���i��E��yc�a������?u:�k5g=���ǀ����`���m���v��7����.2Z�m�E���M�ņ����>h;$`���^'� �tC�L��E-6:\�r;�m�NC�|������,!�~�(��"b��s�����l�����������T�}v�m��Lbp��SvQ;'����]�l�j�h��w5�@b�6C�x�� ���܏���aV"\΁k2C�|H���Ѹby��N�SCiz'��C���Ӻ���  ؃Jӎ��$�mt�	m@��iQeI�/ݍ5���΄뚊]	��B!m�&0�/��P���������dMǉS��?O���BP@��r�w��]�@��9ǻ��BMN}��c���ύg4���<䖆�)���m�Z��P1�'�#���0{tJ0υ@ȅ���}����}c���2i���bwYBlY��`��pr�W;�a��!<�&�d]8'�v��[f��d���iu/��V��ߘ�+���F�����܀���$�.�w�r^��M�+�Fg�q� ��ܾ_��m����χ'I�{2�tce֫��C�f�U��eԁ�h�&��d�8k�	]� ꛻�1�"�6��]�c��E��Yᥘ�/I �NW��W]n����ՠ��!�{�}"��ȋ?>-� �V�a���?j��;h��.��vy������HG5Q�{�!Nf+�u��.�_��D�t��&Tt!`���e�r$6���g����\�HN��D|wT�U��*u ��C�-��ж�>�<�,@k�*���$eo�A{�M��K�/����G�$����F��8zS6f��v��G|��!��懲�&~A�ʘz�N����GׄPL�ٯ8���u&�F� P��+1�O���Z������~�\"=9�\h�}���PG�&T�^��i���?j�x�$܄Mi��I{��p���{�ύ�)��vz�݉K&��(7B�Q�V48�1q�������!�v�Ev�|�!�H`u�Z�H��k�t`���f�<����-���*��2��ǯ#�D	�d;�c���[P�c��EU����]�6!����3l����O��+��<��@����tJz\B+T6k8n�_�lj��� ��;�q��¸��h��jy|� iN�������_=�<�W�*�2/������l]-'d�۶�c� 6����,��\���۽���9/m��ک�[�.��N��#��揪_�j���WA��%���-������cAn��ҷ�� P�L�t<�  ꩎��
4��/�N�b��ѓ�\��8������Ð+{�֓�hp��(�P��%_�X��L�5L���R�]�=K�*k��q�P�a/0�ụ��(��]�Wg��Y�����6��xF�9��AB������ s �vR>�ǚ��g��&`Q�G�`����%�^�\�����~�dh��+��O���~��}�Q���u�!�L
-.�@SNɢ@;ȾG�$��2�a* vp�d)b/1�y&3��0U޷U��"�L�����}K�[����Ȑ���2:�A�_��m匌4���������j@2�K�� V3�mJ����0b�i�Fڿ'j����[�7����C�@̛GJk=�:�p��Қs('� ��.@.Ay��N ��Ϛ@;��]��+ �,	$�ݬ�IPb�v�����Zo��u���1^����Lpvcm���K�8����&�0�L�u���awӆqi��D
�*n��ж�r�������D���Ӆ��t��_�q��O�+��+D ܋)�M~�B�ѽ���QCJ	�W��|�X�R�V)Ne��'2��H�Fj�!1���_�{�>�����c�:y�U�4��z�Q��4@o[�ղ� ��{bW�r�VDv�i:�ؤ������#G������/��9D�l6�:�,�&��re�ɒ�[�a���@�O��)���|���ҵr�RuG����Ӡ��$�������ao����X�=S�{SB����K-���������~��"E�f�����AY���rB}\�a0�D�5��(��?N��wE~pc@�-&�4S���|ca׈��m�*P�a����WVTb�I�]����rG�Ĵ�p����wgD�7���Rc[=6;_�~x h!3`87��,�����m!{4��=�|��S����?ք&�H��JP����aA�����������$Rړ�@�������L�H��qMl(���+��.��U1����?�47�Q>����X���hQ`���B1*d�O>���E�z���a��Q����Mq��_��4�7��b���z��<j�������R5L\����0]��/@-�ŒUY+�VBV��B`��f�{$^�Ŭ��w�2��Q�ؑ�G����A�H�$�jI󾬺\��I�����r��d,���Tx����_�ˮ�*�����#�P�} u*��vM���.��=ѐr�yJ~[T_z����0��G�Ag��S�d�3Tq��h����z�'�=P��6�s.+<�� �R��aEy��] ��ؕ+����,Tv���� J���H�����H�#g/p�+�Pn���>��ґ�E�	5�e�6�Q㮈�6UM(��u����Y���r��Z�y��l��e�w~��j;�o;�����t�iq���Vh�#�tjr\&<@��򜸢�	�R��8 ���b*���s�+�F��J��E��CՇ�M��#4㓫t��l�3�|�l�~R�֏��^4�B	L�Y��2<�2�#g��F�l���c?�bKf��0���lkt����TB�N[݆��~Ȭ�^W�G��3�I�&��v�idyٹ/���<�~�mZ|}r��}U�
�4�v�5�5�i?4�e�����d8�B;�+�&sCc*�s��>��Z^��1�9| ���^�q�����v#L�Qk ��a�Xr:�7q�w:jBW�x�+kUp]�@���{e�-}�A�G��	�ʭq����ol�VE̓�t��gǤ���G�9�㟮�7����8���U�y��v4��ɉJv�z�t���KM�ƍc�z��c�����2#���<�J��|39k�:�y���~65��j"O+F�:�W���h���ק�����R�x-�R����$>>�hR8Q�\^�3�Ɋ����>bB#(��'���ā��1Ǭ�a׌�f��:�M�o-�V���i��
;֬!� ��w����)���e&�ku�Mq�|�0��b'��J��\�U+>��8̳aN��b�?�	4�hr#��2�S�~7��f�x(��Ҵ��{b&ʄ��+��@���*4ۚ9-�Ƨs��O!�XD@G cvMs;�bEE�pPx�oo�[9�vr4�ۇ6�E]�	�}��̫��S�v�
������@���	W	�둩PC5����5E~g�o�Mߜf��v{�?�*�ө1�9�7�i?]���ȵ.|�=,'��~��3md��hگ��a3?Ǖ�t�B%�;*f�a[�T��d�kV)}CCV}�J��]�0V�B��g�7C2p��X@���G8B�T�T�v�+}Lr�,�j}�W�Œ�jv�}&`��Y��=�d'F��c�"���cH�c�4��F�fR���-o85h鳆1�L����.%\mz�4Y˟���������0���8y�p�V�6�G�ߎy�Ux�=gY�U(���.��!*�~c��2,<+C�oMA^�ߚF�hkuj�HCh�1��HۈI�?r�I>��#���0z̹)��ֈC%+|�m�`��I���v���	�D�- ��)��u�d@�K�G��{�LhY2;�@ �)H�i��5o�$��K�}�EA<���4@<�QĹ6s㭑�JV�Ys�Om(��D�>�3���;�n��7�����+o�wr�]���;��Ն&h�/� /J�ٸß��(�s��z��&MN
� ��6_(��9�5�U����������(��1�w�s3�1fT��J7���
;�JY��y�j<�,��*��|��i�w�w�����K����E��,��c�	2�_��}<�/t=�k�W%!V�/���1�̱Oce��zM�6V���R��f%��(���@d@�1[�Ԁ�^Ǒ���>���i��þ�Cxdxfq�^�4�2��x�uapA��k6q�H"a"hKm�TC�K���������V���h��	>EӠ�̰�j��ԛ��.F�L!�$+�+d�����Ut��=s59�@�Y��ʰr��R��5x�Qǭ���m����/Y�~���P��{����!��޽�����mڿ������[�sq�=�jk�w�w�p����pBJ,�ʍ���HR��@��ہl��9!v4� W�D�-�|�{�Żx7ݯ������78W�����.	�=5� �k�4��/��OXR�Ϸ
�]�簠�#TB�7�w��#�0�lOmCe��3�m�P;�����S	�1��NӣM�v$6gX{�d�n������v��]�5��l[���钻���0�z�e��Z(��p�A�0�$���n��3?�r�0б��M}zIqzY����F�ԟFv@�� �N�u+�O�pˣ}hon��|[��+�ؕ�Hw�Q=p�Kσ67+�qk���W���!2��-��ex���"X\�Ec��j;�9�����{&4����|�i0����@��ƿ6˙st����tqL���û�b�����_
9w�+� ���`.%��f�' �J	g����t��q4׬�����㛊���֩�fմ�L8����O��5SMv������7N(��$n�p-�`=SL
n�,;��初d��[-��	:��)s�eA�%��%I�eAo�^ۊ�)/wB�a��̻�b(m%N�#Ń�¨�K���e�9Qy�(?���1��V�걨<=����ڊ{������m�G���c���� ��z+~�X�L���e�D�@�J,�r�������)���e�Ƽw2����#�2@�˼쮒��F0�O>?6p��b�Y���8�]��^��2ŕ��}յUݯIE�Y�����r�s�D0ىl���RIn�'�lRg�[���z�h�~�RY�SP�~��p)�L���`��W��B��:�{�c)>}��H��z[��VK��'Kȋ��e��Z�ɑ*�q�w�zvd�=��=��am��������@WE��hR���yX�?rR\4);��)g���G�P]cs#pG���+�p�����7|��=\|�KM�_8wN�[���H�~R�i�<�����[mV�*َ5���E}}� �m�h����9C��C̐$�m��B��^�	f�\Xs���
{ ߘ��IW���r���t��<S^ľ�q���!�Dޛ ����P\6*� ��EJ6H �k� ;��h�0�<�`4�H�$O5%��~�l��jm�G���S��$fB��:?���#!��K���]�&A؊���o�%�H��1l�Y�m ,�؂@�0�"�bX�n�S8��O1y�B�-��V������"EF�� �'V���U��UE�����Si��V�״Ę�-r���h���mgX�=��ջ	�ȡ�1��=�m6]Wn�δs��7Nd�4�p��X�d�|~�@\�{�_F)���Mr��S��I1B\s?mmP�pQ��<C����<����yU�D�k{W��A��@:x�m��w�9�_{ny�b˵x� ��k-�>�L��vٷ��}$��!)�%>�G|T_��$ɶTϏ-�Ҙ|�8Q����_�$$Zx$����#?��6��%�ȕ��?_*J�xTs�n�E4� �~�B���S���F����>yߕ�k����rc�楸c��$��rG� ����\�;��X�~K�m1�;/�~R�R�F�u��n�M�(w�#mY� EnRG����`:��-�+l����s���a���@�-�!n���%=�M���*���t��7��.(�JҬ���o�p��������y˿;��v)E��2�i�o���
���i�������Vy�w�>�T
��#�T];1 ���Rnv�mS�(}E���~/o�h�S:��=���]�0�
��|^������+7�^�朩2���-�F���mӣ���i��l�<�/�ӷ��Hb�E�Kt��0jv�`����'�'�d�m(� ������S����ؠ�a�6��,b��axC�۵��_c��Zk�C�VAفrf���;!�WɁ�i�l�� �%�{��f\=������A
������3�Un�98�w�bPK�P��iYh�K��P���rU[����2d��a;uS(�6u�x����~&`X��@��R��&C~�+�8>��i�D���Ը;�R4��9�R�@�P��7K&P�;�_�)�?��۰����MS��@����}���G�|t~�7�'d��Pt5v-��VU56�-���_?ߪ"L�*T'	��� 1���bڤ{z�h�²j@���Z�Ʋ�@����!��X|r��lk�|ķ�	%Qy\�� �T�q�OF[�i�Y7�"(��R� �`�ӣ_�:q�`���{�d����3�C�����@�����@\����� ���w@A>�  ���o�W����珜��X�})����Jqޤ���p|O�g��y�y�n.���˄Qp\�E�#�Ǜ��Ï?n��q���ZH ��z���|#d(�UD�����Z�)/���b~��wl�yq_��Z��=�� ����"�K�D��J�X!�H�ƛ�n��*��N=���MV<���Vľ.dܗP��v~�29�Ah�g����9�̥w��ʭ]B��˩.���U���V+������3��ޞ#fƊ|�+3��k�U���#���Ɋ�䧺bG^��GRx/2a&�b���ify$)'��B�*H��r���)P\��F-(b�I��gO�&���n���V��L����������M޻Vk�Q3���7=��vQ�8�C㝋PT�T�&	���C��óx\uE")�]�D ���=�����2\4�&e���.~�@�>~4Y� �x&�%i* ��Rq2�u�^g5&�\ �"D(��15z�U�)�1R1��\[g���� ��� ���h�Q��[*�����;k�^r~�j��c[�� P<�=�"�4��t���\i���F���9��ތI��c�T�`Aۭ=���3tL�6�y�U��0"�5s~`��0�G;�5����W)�����CN�Vj-�vy\�!G��t�Ux�fC�xj5ټ���x旃d�h��g�e ����f��eH����4�~r@�q�+�z�1O�bH�9�@6�� 5��6�WȤ�PF��Yc�m��I�����ݵM�㷏��rM8� �@K�c+k����N+�P�}I�Y�=bv葛i���?u��bi�>Y���@��R�4-���v��-V\��=]l�+��*�Q2�g�� ����~���A�yDI�w���FD��JqH�VJn�9Ǝ�t9W��@��!Gz�a����b�*�U3���!�:Y�HC�jJ&�n��q_\`�A�n�d3,cf�ÐdC���/?NN�C<�r��i.%����B�Κ�D����dt�?��,X�A�^B��d�{���̦���X�yӐ뢨�������3�KR�C��ͥ�����K�r���E�ICO=��b��H��X���[��ő�]���:�_��R�M�.W�΃��:�����7��%��Gƿ�s"{,'�R�k�6��v���"��b��`��L]�`E�Jh�qfg��h�⣁�QhqM�
4ݍ0 R}3_�
ib���"�� P�^ˉ��A���� �B��	�<������b����b��"��XD��o*%
87=�,u��2A���Rx��,vl�;��)\������dQ麈[�g*�/�V_X�p<ѳ<
!��zoMdT̑*��J����� ����, �La�����e��ϸ[93���uڦ�ϸ�,�fA�y �E��޽�w��r5Ѯ($E!��QY�΅̾+����rք�	|�%_������<��/awƯ��^6���:��I�?.<z�1CJ��U1�e�{+4�>���x1|Mռ�U-n��z�hA����`��ǧ|<�;�).	%�u�2��G���&F�g��7�(ֻ�@��B��>`�d2��|\�o:ם�`rc&��z;ߪ��L%Z��"����`8�>mF1?oJ�?�h�J�M���Jj���� Q�a���a����:�(��h_���u�R����us��[�*�o�Z%��ʙ���\6�ٺ��z{V@D'"���Ӹ^yH(��ۙKF^����~Y<�8{���^S$	����mG�S���,?n�5�����w�m6H��s�I��ث�Y��KF����������M�s �84�..�O<=#�����?��s.p� ��(�\�>��Z0y�l�+��!f����QBEm}}�m��#���S��^�3����(:�?�j�Q�	���0�ZN�>1F���p�+���I���uǳC���z1�,���i|�|��a����Ym�ö�oz kP^6ӵտ��ο�������!��1Mܤ1zڋF��E�i��|�)X$��f-��qf�|�U�Nr���nI�Zq}�TBw6�{|y ;�TGi3<�q�|��3�|ڪ������)"#��ҥ���_4�]�A ����槜+z���-�㞯i�W�]�\~W�!?�V.�^�ƴ�n"-�� ���|Ϗ˒G�_j>���d��N�W�3�$<6���t9'�J-+�M �n�$�i�N�T�׭&�fd�x�<�������x�;��0��'����}�3���w*���(ֳ��� �|�"���Kv���txKFγ��+[��V��dh�  �=�S� �Nu�h�YN�l���se���X��U��[�΁V�h�����Z��$�)" ˟$�M$I��@�� �Q�P�������U���A�N)`ie�eV�L��7��Iʣ��Rq#��y�V�M�����z/@�ܐ��%�,�D�N$l�^��F�8��[)��n���N��Ͽ>Rq>{��+`��5B���ho���6%΅�B X�O�:�sX��	g�GF�M,Ŕg�%Gx�6��V	^��`h���~�0�c�����X�[�T�J�0��D��-�,�)��H��S�a� ����&uU���y`���Pk3q@�y'F͔��qSw������~kj�T�""]ŲA�J�Vz��&% �p[��;�A���� �B�B�B(	%����|����Y��d�9֘c��}��1Js�6yq/���tݪ�]�YUPc\ -z.�>������
`��u��Q�6�<�����O��=������!���.�$�4�+�de|_t��V|.M���?G�dX僛����z�����A����YB�{n=kO��ɒ�>3��4�Y<BD}�� 0�Y�
��`�'�X �>��ӒoN��v����p�M�)B������ҵ|�Vog4��G����I�˱~�^S�ԉ��>d�W>���Wll��5^Y��n�fk���FC2Sw}��$�Q�  �,���BS�\(#S�Q�+b�����j���*�~ܶ������A<�)�<֩����}���>� K���0J�2���h���NA晀�z���$8��e��T�N��w���o�QB|��~&�������1� �V�R�HZa�\���˺O�c�8G�=I��8�����=�ݲ_����lK�FɅ&ZkaͼϠ�A @_��Å�n&�gb�V�Y��MdV�+�*U��r-�|�'de�l�BY������4p�~��7���f��|���a������w4��� �����¸ ��@?5��(08pumJr�g�:�^�H��d�3M2s�Vi8��e����oH�Z_��;x��h�?��vf�X������U���֣�c#�����+� �)i&�zO`�K#Tfw�����w.���O=&�n�f
�Q1t����A�-:6�ED�Q�9k��]�\[}�Z����&E��L�IY0�����5%rs{���*�.����;en�hm����7a�i��H]I���(_��In8�f5��Q&p:��Z�x
i���֖���pJ�S/G��Z/�9F��됰�}h�EE��"�;�>Yk�w}�@�a�r�xy�x:���[�5o��B���Os����� c�+_�V�q�_��xN�|Rt~�ss�焣����s���ER(�4��� ��} .�"�=H��޸��'���M������]�Nêy�Ẩ�?�=4�����Xc��f;7���r8.D�R�dBr�L?T̉p=�����Rf������l�o��l���俒y�fG��M 1Jf{M�� {,�Η5�@Ң��w�d��#۝���Ek)q����w��X�����I'�C@����IF���Ǽf� ӕ~dԕt�'̿������p���|Ma;�f����EȚ<_ &f�� ��Ar������o��|w�����\��ys��<CG��B@IɅƘ(P�*b�� �}.�Q��%��ƽn��ýj��An����=%��眹��si��]�~TĘ���@ׇ{pu�z@$�{W�<��?_��V�j{3	���쌕ݱ��#%#t��9�uOۥ��!qi@����Ԥwq���ʛ�0�,�}@V-|׌s��M��A�a�����Q���iY��Q�UuuU��8Y��@�,���)���ar��e�M���N��ޥf�+��K��"�ejJ���������,��E o}������o�IDm/�s�D���wJG����- ).�%B���ֆ@~�m-�6�����U�?^�*G����������N�Ƌ�؈Sn���Հ��}����F��6P:Y��ɠ�% S�g v��.? N��r�W*a���P�Ep�J?B�A�`��&��l#���������Ğr�*� ZY[xܲ�^mJFD�^����-��sW�2�����l0қ��g[|u���^�G	~m������7R�$sF��E��VE2�Ҁ  w ��ʳC��	Wc�C/%s;G�b�B��FR6Su_��,� e�5��CM�P���i�U[���K�Ү��+�&f����	�i�b���j����%H�@��B�'4i]��GQ�6�Z��� ��7�`�������P�d�B �	��" �������2��Z����l_F��k�j��ir�GX���r⓻���� �d)6m8��]��(���t�����Bq����p�#"�;�N�����E� ��Bq:HZ$��,����?�~��!y���mk����J˧�0:�T�ŭ�n���D/o/4!�Zu�/��w��셅���hO�C��Eܔ7˱����N�R���+������c��/������~Q�1nH��m�,��l}��[��F`�F&��+�>Q�����A��c8�rf�2��8�q�Y����C,�@����_�����A֣	��:�#(��w����?�ghu�dV�&i��͜��
{}{m䚉$.��J�^Ib/,��=&�v���!��6�t�dO/��j��Էo�y�������35��jYb�ן,.�m�،SƢ]cB��k|0W���ZhtG�e'٢6WOArz׽k��4��MW�r��u�����*�u�s�+,�vz�	\a�+��7.M��2��q@�N2�e,�P	�	}�2�#"F0:�̔�7Pl�O�8X��c��U��ڝ�wb��K�h��6���c����}͈� ���C:�@���?n�(�W�-W'�O�t���YX��֞����F����غ
�� �\1N�x@Sڃ��Nh�nq�*�!(�a�[Pa��<+qF�`Go���nq�"�;ɟdH�e2P"@�5��H45;�j����z�����w��w���nw:@�RF����C �{ok����D�vSX�]=�B�H���v���2AL������%�	C��,��#^���w��f��^��펋8 z���л��J?���ע�S����H�+ɧ�b��g!��`�ѯY�Ε\֍W���~�R�|8���)��K�#�N����p��%��H��:N�U+(kR�o	��޺ͬ`��.���ހ�����h�ngzȣS'sH�-�5��vF��M|	sw�h��o+�-7�F��c�4� �?>�>����4���U�����^+�5��KF��C(Z8W��u�x��`�r�B�i,�U�+���.A;���|4\xO2�c݃ۻ��?�/�YCk���mY�T�v�B�]B�jd��8��T}m��9��?"�I�D�m>r��^x���	,Y\�m��ח>-՗���E4Z�8X<f���BZ$f��C9"j���CI�'�o���L���������'��¸�׈Q֢<7���(�_Aw2�����!�kP>�+�7b5�����b����s�j�Xnθɗ��2��U(_e��qS�B::�h��p�māۤ��9�n�{zEn!y/�݊�����^?U�D�W�X��"��z`F�*�0�U�5�3�����3�!*��ũ���[�ei�
��q��3A-� ��"b]Q]J��rΥ�UV�Zȍ&��|)Z"U��|dhi.�}h��^r
�K��@�Vcc�Зe٨�_� #P'�A@���=�a�5#���g��
s0�@��,g�NG���b�eQ���li�ɱD��¤��@��%����zn\/�:�����#%ˋSH�o
�t������?#V�	�{#�X|�Y˥�l�޼S���'�f���!��6��Q�,R1R�Xn~fb����ML��Um��%�|t��
���Y\��]&�Ri�����ǘJ�����VV������� �5����s6����PL�z�	Gs'fӭ���䰊F!bO�F��AXa������9�O�}���d������W8���K)��7Z�����߻6���-�%�����X5�?N-Է{Q4:�>ҾfV�97�5�V�����zK�Z��mH�)���!��LKf�n��J�M,�MI�������e��aܾ�A���U�=���'��V��":�76e�]��v�z��>���P�'qT��5��ک�q���=���ܓ#��'Y�ů��k��`C��F��*�뾩��n7�f�R*AO�^��i�e�X}��>>(4�G�u���s���T�ɴ�NV���3�n_X�^1}2=̫/�V][��.�'��T"�x���p���� <��M� ���]�F�ur�ٓ����������O��S���f����{�W�zd��e�)\��Z$�KU����V+�ܿk��v�?�ܩ	��)
�AI妆���H�r�h�N]Ӏ�LTe|��'���j��*U��	5�qO���6� ��w��H"!Yll<f���/�c~f_�����Bn�ŪG.�����
%������wN4�5h�&�3�����Y>;�dnc�4��x��/5�+Ne��\nD�2��; �5 �"m�I�!�����X�܌�#�9KB��hZ&����m����$�e��v1�Ū�9������Q��w �ѕ�ܐj��S�����X�`^�#u�S����%3���h+	������,/�7���U�"	�eV>7��p�9[m�r��e9��Im7�O�c�F���,�=�ѳ_���{����d���n"��`Vv%� 9b�0GV��=ǒ���KyNYI�n�Qq���1��wZ����U1�.[�q���*Qgb �0���c�xHX�Dͫ`�׿T��
=&�h���WzP��!�:�r����z�G�|0�#���k��Yb���|
=�Sz
�	���9
���.�m�)��L�$|�rz~O[��$�M�ќD�|�ԍ��m&+�k�d]'�����r�\���y�Z���h]þm���o�Xl����5�P�c����S 7W�{B�,�
������4{��-�.�,�U��և�l�������Џl�~)��?�J��=٭̐eV8�ɥ\G5�ݎ��-������Yڅ�5�p��Ԩ_���	�8��).���O�%�%�0j�|wf�r�=����3��0��!�D�q�~�8�:4�gJٚ_���͜q@��dnKV������]d���S�r~�l�xs���Փ{9����~/��{7���y)�kO��Z]<a��Ȕ�%�O8���Mi��$U�o%��G}�ݖ��o�	L��G�[���\��D̟�	�q1��N��4/�U8R��P������X�ɛ�#�|����������vS{Crظ��g�n�dj�Fσ�2�k�ػ>�����6���کEϖ:��-HWDS��V�O�z9j����Z���?�-�[-�L��N>�ܻw傦sA���!+O�?�B�/,mo�������]5��)�fJȡ�e1��e)�ܩ	(ٞ�"��3���빖��B i@0vx�_��$oV1��#om��+R���#>g����)A���Zk�y�_�'��G ��J�D����YU�����4��y�y��C`ɪ9�'�n0���,eZW����o��7x�+|�������Ig��'����%��B/W �07!��?fWW�8�PT��/��}�<Se��g [>H��؆w�(R�ɨ�����g�7�e=�R���.X�z���b��$�(MFE�)��JIu/��h�{{ P|������K	>���ɇ2��㬺s�{;y�����'|���+�{�n�*\ǃ�x�5��n-�h~mxՄ�O�?�<�� �����Q��sE�"FN}���U&��ɓۂ1@٭8��}�g�=�8����_u�9|�Z�A�	S��cJx�9"�)Ã�>�|�J4���|_�������]����S`���t
"5�)z��*c[�B�D�]K��I�q��HͶ�O	�2���Y��;JYU��HQ�}]{�&~�Ē�Ϗ��~d�L�x��壂o,�8!��,��^�t�tX�FY]�7������*ųa��$?ق+�ߟ��<eF�rmm]����]�߭�0�SKL�t�J�}nHX��EU�.Ü{ ���a�5�R�~bq;^ ���Ğ@{G�Ը�T1���Y�dݏYv����: _*�ճm�M�{:���۔�-gr��ҋ�c��Z�����@ $��s���z0D<�1���q^��f�����C����P�J�<�3�����$�km)a~SD�-v!ح�k��Eڢ�O��¿�/AnQ��GV�9v�b�,
��$���lf� �=��P�}X�� 4�0��D8-sƺg�D�S�m9v�PR�f*�9��
TV� �!փ]@*l(*��,%�j����Ȩת�#�aG#kO ��B��Rꮀь���Gk{l�_o��ʦ�)r��`y]5���������P_�{�曙b�7U:f��z@9h��mG ���RFNA
�� '?�:��]�w��}o\�a+�k�N$���z���in �@�;�����e���%xS�.�1"sGơ?�X���j���ژ@ρD����P!���2��u�K,����e2 ?���B|������aM(�V��R��kG�{l��ۿ�
�>��p3vqؤ�f����z6�	���6�\v�k5a�a�y-��G�:Ŀf�+f�]�)r�x�=���ْA��£��ʎ'5�����~E����Zl��J�L@ |�����r�>�<6I��P��>�T�a'Q����ۨC�<��{��>�=��y��V�
�!uw��0�VD}�+�:m��j��mtF�n��3Ĭ�h�֜���=����5Dݶ9��c��n���c�1�{2c� ��6���B6��9���T�ᦱ����5H�S[xَ�$/�zK��yoz�p�l�@�'l!q� �t�G&��Zl��&�����X��uM������<����L/��I����Z�ה>+��45KG96ʽ9�y�Z�A/�.�j8q)ጡD�rGȆgFHuYk��`=xD�9ҏ�&�(|�h� B `�T,LNPd�D�r=��V�7���-�n��z�oN��sY�E>���`?n�`Z�{�+k��[�2�/�A*�  ��I-�24}s03h�bm!�ٲFG_��T�`f��˟y��~��5�I���� ��|ʃs����1�Ky���F��,��!��)�
ݨ�88�/��](m�f�&q��fZ�� Pn^+��LD�bhƷM�[����6fC7;������#�+( ��8�7��r�0o�*0AY��Ӛ]IG��B��i?7|b�L�WS4�o=��S���.�xct�U`y�c?���������V�"Cط&�fQ��P��F����H¾ v�� �w��fM�ܣ��x,����"��}AC3�&Ӛvt�ƺ�3^�|H�d��]5��Yp��v�(�˫��
�"�b��[��B���=l�ލN�y�k{�|�:,R�j���a�� �}���=�Jh��.�"�dgY��n���o�#}sx<�����j�Х�ڻ�^ �j7d���#"�F�W��e�(�@��D�� �L�y,J��mnT�Ĕ��;&ԷS�c�#�np-������$�
��>�(�p��O�BЬ�2�p�%�M�j��R���Om�-G6.�L��<� .۸�՛�x(�g��v���0=���bFL�i\:���N��KBk���1�%x���E�@m�-K~�a����py�=���z�x�y���_��y6�
��P��YULݍTpڛ�]t��'�_L���o��]�t<٬R���6��M>"�0uU�xX�9�#W8���ݗJ�����������k}*�`�������3e��f4!p]�N"��zEB�߹���;�A|?�v9�!l7���HP)��8�Ӫ`~�3�	fk���`W�����!���u�L4��#(����+
�cQ�2U�t��	��(Y]�����^~,ع#��ΐ�O֍����X��H�v�X�sE��D���:������4�'���]��
7���,��,���R&F������t}�e#��q�pь0"c$�}Ce=q�#��n��El�$	�>��,��Cy[��N���_��.-�$H��F�A����5��]!���XM�����U�;ou������5i#VjC�vT/ݑ�ss�h�vC�)S�׀����c�q�8!c�����G�϶��G�w(�vL<:�#eC ͦ��S?���mLȢ�<n�lc���)�y\j�@�t�-�XI��j��?'��:�x�I��gi��\d�:Gm�h�hN��P����Џt�v������")�n�X��\ވ�<y1b�4=lQʮ8|Q��p!�4��{�U]��� ՆkhL![L�*���0���#V��?��
�8�
Ůjd���w�k�=������-O��ƝKqN�7z���T��$����X4������%��E�����v`���9�hB_�#�2�����<�=C-zcR��������T�b��2�y���z�#s��]C_K܆7��N_����/%*Z���t
~r��9b��g(/�(vϒ�<z	��ш�Ͷ�����&��H��ܣ�"ћ���%�_Z�z�0L�����eɑw��+��|�O"TyE�t�����j��������U�u��n�}d��þI����)Q�^.�q���8k�}_�/$n��	0!�T�(G��îl Wdk<��u/Nm{r~��Z&�� �� G;$n5)��Ӑ�x��n0�aO��r���s����-�\���v�Hҿ74&�[2B'_�һ
�Ý�r�S�[��9K/�ras��Q���"�K"�"`s	�M�sO����Y�}H�����Y��@~����0�1��GX��櫶�M��"�d$س� ��۪�KF��b�v�y
kM��ɽ,[�_]b�M+��;���( -	_�<^�ur�L��w�C{[��ʠ�ף�������2^c="VN�m1��3B�:��@r��-��D��־����§/X�m%-��wf�v+%��U�
h�=�;�P��C��/��lm��sզ����N�؅h�Y)�Z��3�8���?-y|e�
�F~�hڨl��`��$��!��7~v�@@����Yn6,�{鳵4ҊW����N��oF)t�%f�K���������Ҳ�V�B{a�MM�$���֖>�g�+��{��3�0U�v���-d/�gȴ�h�(�"����2%�>&&��{��ieϖRe�5Y���2����oK�j�<5�W(m�6��\���d\��ª�������yO��+��N�+�o�;��'C×��q�xk }�"n����l{3�� ��l���/º�P�S�P��+����p���2�D�<�����L����~s���j�����k]�!��ss����V�$�$���`/��;bΖo�"(8˭�@ժnfwT~�=f���q�2�8%��Ĩ�`��S��ޛ�o�,z��:�%씤�d������x~R�q�������?;]/��O~��<�t�ťM�94�T�Uj>�hm�?��ڍ��'W�o����d�wj��܎�c*�й�F��w���ik����(K<zhf:έ�0�&M\�dǆ�gee�9#���Rp;��K���p��8��i �Z�ɚ���qV����w	*)Sg8���Z��fz���A��7��L��^�U<<x8����Uc�TВ\7���;:2&�tgɢ�1���u12��;(��F�M�B��]���D����Y�V�Ա�݀T�FoqX���UvɫU�m+'�r|?�l����֊�ӯʗ���b�R�Sf�>rn�Qe�cv�]�'Qc~L���wBp�z��?�a{���ą�C\����f{��ODl�o��-JF�⚫��`��R�{��"�Leޑ��ʨX�����JI��b\�'�1K�̚2Gh�l���]���>�/�J�Y�ro0[o�y�?*q���Ybq�(�n�GZ\RV��QE�g�E!�M�LuE�:�����g:��"y�����'�V�jDJD���Sl�/��J��^��+i.}:RfPC	%�k�x)�Ʋk�"���޲�WkU;ܗ�s$KD��+V��G>�i?�z��hI�����PLr<l�Y�� >���O�/��3|I�k��<a�K�K]oTZo
P	���P�2\�Ʈ�%j�A�� _�=b,L�:�l
t-Y�ֿ-�0�݌q���؍��ͳS�?�i���E��݆�Ss�OR�&d�Ӭ��Ȕ��H���^��q�|�ĝ��+���8�~ɩ�r7nu�I�2�f�%bv����5���ٞ��^}�w��6P�A1�bmJ�/C�xh�A��	�R���'n�uv�g^ Gj��-��YO7Bk����"Ib�+`�c,!2Hs���� -=�%eα{��s�V��<��N&g?L�b��`�H��;ܾh�n��[ǰ���g�D?B	{�;!=�hEO�CH���Moh`q��o4w�s��^;�{���%������L�Y�6�h`�^]h}<�B=����d'ʶ�A�+E�[eiI+b�d+��3�{<4����
r��!{�������\���'6郋��{�v�m��Yj2i�+�L��.�V�K�4���|/�f�PV4/*IBkzgx�v���y��]=��^���5��YuU��|V���X�{x�@:[��)Nр������/�~�\:$Դ�Ȭ�P�}C�9!�Q��Yl�OC�7�U��Z��3��*a2wP;1l�K�H�������A 5�eá���0|������2�.@^�zy�%u9;Gǯ�ѸCu��Y�q��j��a]�1��w;�Z���6]+my87���t��>��ǣ�:�ƹ�}�Aq8	˯�[A�6�S���ˎo�8�:��:����Y.�ȶ9j��~�ӊ��o !�g�����T�A�
��?u~�鋜i�r�՜��v�hs-&_��]��@{H���j׹���v[W'�̲�EƼ��F��r*��̱�K�D�䳭qIS��3�z6�lє�-�/)��A�3�M�C�.�7����^�ne��L�`����et�������B�U#`h��YT]=�h���]y��)�I�U^�#�=�r~�Af_4�y������`�^����'���$0�\_������c-V��${�U�����j�#��ʳ��	��~G�,D?u�y-�v�M���l�G�m�3F��ٺہ���h<��6����kak
R����FwZ��r�%Q�cc柽�����n�*��N�scjss�ڋ7�S�Bef���O,w�"N����������m2��{I�
A�?�D�AL"��d o��L����v��!5pS��hi��8��k�FkĐPO�rW2H$���vg����(���izrKƂ�����MB}	�5XN9���G�ì]�-CTH��Z�w��*�Q���T�:w#�%/�j�9���v�Q�I�������tb�|��S_��H�6h��ܷ���z=EZl�;:��$)����u���[�M�� 
We}���3�K�A�p֑�ok��$�!�b4'�2?�=�Q�3�#��?��΄��ys|����9�[�����pjI�xy�v�{��C����|�T�Y�s+��Aހ/��9ʿ�+N=ni9�Q燈����I.)G���ӊ�<�o��ˮN�A�Ƣ����-�����3!W����QP8���H%X��yك`�\�!�)�J�P����Ow~i�G���o�7Jw�G���~f����|�K#��9x�_��oS[+7�H��3�{�fdZ|]�^�.h��5�St���2u ��S�ӊy~�^: d�CD�ɭ��/؃)��[U���:H�����+�=n�լ���_"�]ב�A�1�d+�x3�����z�/�b���H�O{�J�ʧe���]*H��9
��A�Z�����*�b'��xB���T���������JFߦls2Pg���4���-��hKM��i����Ґ�Y���(��2@D8TNS�K��h��Zq_�)�ҍ�TL�Q���^�rc�@���cW (Ms���r��{+?h�J4��s]� 8}X98n%{  ��E�σ"�Hu7�W�wL����F��B^ԭ}���A�)����/4t>)�[������
�U�]u�`#��&""X	�橴�'�D'����(��h  ��YM�
e��Jr;�ہ8o�K�o��Dw� �ǅ_���{՘j��A|ٲD$�<�)��\�~xd��|�I_q�ҕ��$��̡���o-�x�:���{�A�¯q�[� �o`��%1��]z�F+�����dI�#ɫx�G�o�������%2Ҏ��e�^� S�����CI!�} �g֗ߟ��N}��~���,�~<�|�ko*S׀jED�BL�I�?�Ɵ�� [�#ԎYT&��^XM��HPi��$��&T������j7�X�����o�K�$�,��R�-���������|�6�����3�Y��;
�Fv��G���s�U��>#ҫ��
�:���Ď�A�K�Q��3 �ĬK��S
�x�iMw�0�$���$�v �!�Է��U��B��p�^5�6�����[���+૙������u_l�}��7=�����_h��7t�}�]�������A�4H���>����n�F���#ɴ�1�GP[�b��l�Q�9���rlF�%�wJ�[J:�FQ�K��6l��`���$U���D�"�ͽ;ֹ٘�AW����I�]�PB�+���
%���y��Q+��H
Z���3�_���(+W>퍨�­�K��FN���J2q�䭰�u�{e��A�I�_����[�E��.f|�=�b'[�*��Qn�c��ϋ �CF�5K�9`�����mGVR�\V��K�/(�B����F��f��M���}疏r�U���^���v�K05�����0�8�v= ��!��!^�"�B�N}��WZw�~y��ᵹ� ���胧�Wk�]/V�y��#�����'H5-��l��ytps�m�ը7��������L}��?Z6�,��YR1V9�ȥ��]��nY�4'l#N�3��S%�s����z� �YT���d�y3[�[��;�����[��}m���_���땗m	�㞟B)Z����.���-����ރ�Zl7�7�?$dU1��;�
�}G��D,����1��f��=�=��o7d���J�����2�;N���	A_��?��ͳ�Q��9�|�l ������A�ŋpG5p췤�m�y���]�Ŝ���G���m�㠛��Z��q���+�u��j����7O�����"��ٜ�w5��*�m��\�$�Q>��
��]��Ɵ���%"��Q����m���v��J��R�>�w������W��}���Q"D��`�P���[�d�|��
��6dЗ��XG�n�Gv���8?���ȕ0����qAA���ޔ�a_�4�UWߎSO�=��y�!y�O��S>xܩh����:���`�R���iT��+�W����}��^��g{#���ݢ�'�Wqn>u�;���[��y;+B
�屼�W#D=o��h���1���rW��e?ﰐ-�䣑Bo�C!����>F4���'�C�D�#��T�
����j;O=����$�|K��"9�'�7�<-wx���u�Cˢ��L�8Z�M~}���+#�;���p}����Z7B�^��qk�U�:�UiZ�A�E�]ٿ�/k�ow�8R��Pk�k[�{&��&֍0U�f=U�_͢�)�k.�T�*�*Aq���ُaSZ(��=�'JM�+�!�}^�JB�$��j�9��[�F�2�,��;����z�.��E*\ڜ��kc�����/��d�O6ށ7�UM�tt6bC�v�ҍ5��^����c�$6ń����h�9�������lV�#�VåS&�oϢ	�I_���0>o��Eo��+Vސ��`�2�8��.\ƍ�o���Bh�
�+������WR�#%'�(���a~��P��ܺ�٨��h��_k@<k����;.�nMw��d=l�ӧ�ګ�W��������k���t9�ԕ��{�5]�_{�q �^8�)2k;W��U��&�Uz��Yq�W�A������a���
�O#�`���$L�_��|��Je�4h�S
���.*��1�����Tx�pi�Q�)��V�6�.1]����m�Ϩu�V�l�^O*�v����Gk#0%��[׮�(�;�dB�"���޷z����R)��*��h9R�����~}F�9�c3��`jw"�����˕c���������J��)1g��[sxd��~lg	t�p�O���@*=FQQ@.|NLw�a���{�4��Ny~(9��x�A���"���\��a��u���mu��О��l���?IԸ�ȱ����h�-�OV)M@�t=�������ҷ�Ny�ZU
5�i�,��O<s� H�>WS�Z��&�S��)Õ�zn��E�]���t�C
�i3����Z�^y�������\��6��v��5����.�V]I9M��5�Yzu�0��Z���IYK������K��+�N��K�~!I��'�I7�ɦ[�=4�-?J��*/���N���oe�]����J�9դ��l|� �nm����K\�ғ�q�r����Sj$��fD/6�C�f�Vi��7y�H"��x�r��LvH��v��3���[=���g�OH ��5H-�2�����2צ�e����L�>'�seId^ �H~�N�B�{�*��ǥ�,rD��e?�I!������6c�_�r��tD��=rm^��Q�,��7*��/sg�
�N=+�1�B��%y=ZԖ����N��ڮ|�C �ݯst��,{39,���]�?�Pk�*PJV�{��'�'k[Wi�8#�M��gۋX�-�[RC%���g�^�"�{@Aq��t���=OT&:���U؍��nG%E��f� !%��:�Y@�N�i\yt����y,���u�k��~!�ɦ��=[땝S��ĵT?��%I7�/��+�4Z��G$R��x���3+���� ��1S���!�aA������F;e% ś�3��e���]�<��R�,K�v���`a�`��ȷ�/5�y�j��0�i�
��8�*c�fK�����	���G��=��N#^>�
\�o�Y������b짯��B�C��J�y�D�h�5=���oQw��Z��WL���ݔ��n0FTd��mgLĳ�]zQ0f��JH�7�TGAK�J�����K�Kޱ=���Ws�p��r��=jj�y�����s_Z�[�R��>���\f������>���V����sU�U��#%��v�Oȟ7�jF�o���{F�z�Ĵ�|��4��:��X�H�����3H�������'MO�[2F��kU,�S.*:h'���Z9�g$o,b�{���$��a��%ݟ�ť����Y�`��<Yw� J�G�g��9����A�\�HV�H7(5G�4�S�O��eld��vb`���=�՛Ju�$m��R�И�_��扽�-p-���gȶ�G�Ol�WP��Q��N��A�Λ�7Y.-�Z����qIq�;���o1�XaBm�6xw&8H� <#��tMJ�@����&�*ߺ��Q��N�5�*��_�{�� \��S��sp��)�9Zi����^���@���1��h���h]!5F͖=���A�;כ\C퇚�U&��?�����,����[]��%�ڭ%�Z�^8�O����5�Y��8���y�b�/��/���MW��ʵ��b%�o���Lci�[�Xc����W���z�X����y��R��_��Ȏ0Ս}]h�˨��˨X��Ս���{<Y�� J8⩊�aCBgAA���gzp�R���5�lg���)ֲeZ �W��DrYQ�<�Υ:��\���˖W#[�������/�Ϫ�u�j}���n�43�������V&l�j�So�l��:RΑ�˱��Hx����5O����v{K��u��W�O��$Y���K�ϯ��`X:��� .+K؈|����e��l�ʓ�wJ�x��uˬgoݧ��E�y+d*��:��Y���E�߆=J�.gd��⢘�$�*�*)_n��=R̓��,�Wb\�.0�h:��i�bϐIj�K�*�/,M�����D�>���&�eI�ܜ�����S��!Oc��;T�:��pB�<���|�MH���1/dj�&�[��R�4��0Ex��:�����V���� ��M���`�X�{��O�3�拆qZ�[��v.'�Nж�`�XT�����b���s`PP�ʛ���[=�~�	���f��9\fcZ�6�u��d e~�6rS͡Y���j�����i:�%��K��'FĆHޙ3�.[�b�"5�o#����I�I��G<��Wp���N��^9���1k�;܎JW��������c٨7�[�+*��R�y\�W|\7 �t�D�hR�6�Zzyy���9�O����{ua[�+$��h�p�:�$��W�:rk ��#6w���> b��y^�xYE�����kjj"a�[����t=)����8���e�ֳk��'K�y��U�S)�N!!V�d�/���g�&�f2xu��o9��n���{���v� ����Px�����r��&�%�%���WD��w�M����ګ��I;��S��
%,�J˱�C����ޜ�|���LO�}_Xߺ�)�/^�������%�ѱ�����'A�>���'�a_��yL]����)ݩ[Y�h��Lփ'���-=�SMS
���g�,1��X�l ���N/��M5�5�o|�-}
��V㟅3��̴DXx5<B�qwRڬ�[�L��Ŗ��o��y:}��
Њeku�*o�ʵ$�^8�+�Qg��L;�h��o�b�#��F(���q��������G�±�ݰ���������L7�v ��'���v�B������B]ϰ���%����Z͑���+��b�9åBI8���4��- cV��u <Ƅ3�B8O��w��-�H�v�`1vk޶�_�����V�_���
�V�ZUo_���6���}����h�7GtIq�r��
 B�˓�a�L��zc�[~냤��P�9�%�w���Ѿa�BIk:�~_��������WwW���(!�W3���W/����b`�V=U���dV�Rq���{/�h���b!�jA������aڇAJI�n�i����EJ@J�n�F�����\`	�^�;����s?����{b暙kj9��ߡ�al��Ѐ�OM��� ��&��ޜ�As�W)h���z@z��uD�t�5���ZT�3��e_�\v�'�
��9�JNϸKV�F�\cK�/�.(O�����"#%U��1쁱������0C{�Ɂ�,�J1iIv���/� ��*B��?�@�;�̝�g.�'��J���xR�2�7q��D:ﻶ�l���z{{	��j���"��b0|[r$
���Zu��mP.�g%w'�H��xl�
�̔���~L) j?4�l������}���N��}�˧�z�%?!��b,�LJ�)�k+�f:�O��D@�h��ϓ��ɿ_^��x?;Ѻ*�0l`&�8ɀ��~��@Iɾ�����:��YN]S�r���Y��{�Y���?m��-g݉��<�S�$����dZ 3����$w��˖��/��F����۔rB�܂�����f�<�1d����+8�`��G"1���<�:�7�{K�=�*ǥ���C��ؽj�/�A��l�!,�km�N�z���u��ܪ�1:8��Un]��e��<"���Ĩ��	��]\]��vJ�IQd�Z!Ȓi[;��,�_�:���������\5��q�E!�9W`�$��s�+g�󶅍���b���*G/�X�{tAY��>qO�i�jz�w�I��g�W�>��ѓ����MČ��.l�!_��	�hy���b�	6�1#X����Y��۝���|�z;�/w��s��� �Su|�@L@��^懃`��R�"��诶�o�Xl�'�V�K���-u\�	��]��=Ri����t~: F����@q����5"���;u�}�)lJ��16W&�.X<O^�i?�Ѧ��	~b��L��!D8J���Z�wu}����%&�W�ޞ��j�/7�^���1	����^��esj��n���f����T�-%c�q
��:״�m��J�ڝ�Z����L�z#Q���\ʧ[vk �MAL�@�M
�M>۲��w�5h�y�8���7�<����#�Ib�d�FG�]Ӷ����ֆ��|����rߧ5�1�̨J6�^�����Y�W*͒ADL�&��ӯ��3�+ \��J�uC����Z�yE�E��1��0D��05�����Wy�������7ָ��mgNBe再5�S��Z�	q�G��L�W�Q�����d���*�ɈS7�=�C���Q�pc����:9Ū��gh���W�8�hg*	U�ۊ���j\%Ҥ5� \��
"\R��u�O�烷i?�)��Q�O;*�mn'�a�3rTx��:�Q�����mZi���O���j0X���J�lJ�Ze� �й	4Ow{�Dd��a8uىA��V�jYK�rM�֦ٵrn�Oi�V���׳Krr��Z>�R���g�u�Ũ{<�drՍ��O�S��5]W�%0�mؽ�"�%��%aGwD7���/�'��U���1�V�(^��S~�jC8M3��v5�`�ș�W� vG���{�u�_BA/�d�}o��>Tk��UL;���r�M���Ɠ��,�߁����#ʘF���+�O�"��A?-�\�f��*��'K+���&�˿���db-uCW�����Z^B$�0�m�^�P�&�遡Ǔ���a�<��V�x���G5	���ұ�<�ê��b����]��~*=lk4�d�>�dH�~Ci>��!��x��s��|�K�e�'�5��7�8��k������R�s�4wY�ym�s/&��)%7w�3 �)�%��"%r�T!��de{�U�ggB;�x}���!f-,,���g��H�H�"m���]�QZ�e��SC��zW�,�_6�ô="��fg��+d����P=����8�����l��HJw6]II)#��'k&���4�x%��ꦨ�dL^�|~ue���1b1XT�5�6L�#��H��|>Q`�4�G��Y��;��s�)z�~ɹ��]��:�r�eC�f�P�>$�;*�o�.q[�TCFQF���'q�p`@��߿^q�ǿi��++�N��kJ�4�F>no�ʙ����u�_�\�2��O@@Vh9C����/OP��4n�Y#��&MĎ(�i�@Elv�! �G��U.\[A�o���/�?8[��}��5 2;S�V���:�++2���^���ج�B��먍G������ڧ�V��`�\�4������<J�ի>�Ð��֡Bq�Pk\��5 ��>��E���(�*(�aйP��݂߈
`��|�X�y�Ix�g�i�iو]�P.�-�E�3����_�ܡ�33��?$p��<��j�gz�j������FX�]��j�\����y�X1l��0c��$X�S�x���_�e(��N��c�ל�Y-�#/���$z\h��c�Rա"�)����vNN�2�,ƾ��Oy�'Ri�Z��@D|u^.=��AD�A��S/1��v�_\GW�"ZIC�'&�+4����zx�͹�@��ڨp u�]ܗ���l�6�k�v��!��%���h+///>nۇ�����ٷ���e#�Tb#,5�,5���HST�<\�5joI(K�נ�n�8�#��ҢSWsA��Bx��>̛C�ɕ5k�Sl)��d(;x<d�CY0����klt��^̬.�k��
4o[ӤyK�"TvZ!��$��ӝ-[}��!��p����P�1gu`�!>�.��kohP��7t�����zآDݶ��B��VH^K�l�1I�w�L�������nd+�V�D��6+a�b���@�Yȡ���\	����R��`tO�׾!�}�bk���U�䫬�C�4��;S�d�����5I�?-����+��3��%�vy���:�9�]qS��(:���d�q޸ĝu �6/�1�1@߷朠� LgK�Mle���8����F]KG���6��(:��<)��K0HY��ϴ�������L�OB0'��ب�Ӻ'^gߪ�_-�D�� �3QT�zI����m5&f��(��X:A\"����H��Mw���d��Y��4����7�V����?���m��J����95�|�a	s{:���Y�k��f�5��C��y��	c��㶫g��b�5�'=�'mW�̟J+$_����OS8:8`H�g'��Xs�1�_ܑ�ގ�778:t��ϟ
X�
���z���Ϸ���$���3�~�z��U��y�{Z��߯ɅO�jm�-@�ԇ4h���E�M_��9�����,�"��C��������n�s=��R��D����f���Y>]`�����QM�i����>��d��R

-��cI^���/������r�V	������2�����dLߥB��w�)djz�oi����ġ���<@s���*mMw�U?%��6ߘ�uS>hq:2���C�x
�Jk�Zl����^����r��m��`#	

:�H(���!.�;���q|
�Q�1�$��]�{琽��7���K�㛪�1C!��O�)�p��\c�B�� �G��N�2Ͷ�S�����ǟߎM�DȬ�ܫ d#~���T;� �?ň|�X=%��T�/}��m�|�1���7.e,����W���U����'�edP�����c�kq�LuuIB+���kl��0���]T���&=I�|kּ'���c��M�v�ti���HHHzC'+�-��oW�-(��/��1B��A3E���2����X=�nֶL�Ϯ�4p직� ~�W?5�'�`��%:P����s>2J���UT����������j��/ *��k���&��!p�#���#k��
��efŦJ�R._�7_OG���뫄B�x��Lܲ�kQ_!�\��e)(�䪨�V���M]�-`eN3G�Y��5u�P�]U����O\�������|��|�V����{��.�ټ�dJo��C���*s ��`��D��V&��['.n�7�2ك���?Tm^�;R���)hA��6�>�r'��/Mk�ī_,yn�m_��(��6�pf�D�^>c���M1&p;�%����J$DEB:~�k"�u��w�pKj��������|�����.Z�I����8�
�qx�r���M��dB�D,	^%j�6$-9\=� @Z��=�zK�R�5������yS��Lx�p?џ�Y�x���JWݎ�yO�Q���࡮� """��(Bj���U8�����.8��1�܀8�n��� e�_��)
�<�����;�����q%�	��n)��pϧ%�kƯiL��b�.�ap�_�'#mqr=T������x����0�?�^��v3&ᝡR8�H�U����vvl&+:�ְ�kDQ+�+<_+�
����������Ÿ�YD�&2zt�&��=������y���
h҇�w-2��Y��e��$�-����6��FYx:A��</�0=��U.A?�K��䢇�̳��q�5�dۮ��{'L��-�-�[ڌ��.�U�fg�m��+���,������N�ŵ�/>bh�����<�XA��֝���~[�(�e��{��x�r?�5�ֻ?�`�H3�i�U����iZm����"Ά즤��W[C��gro��k�q���J������S�R�3�����-���2c���3Pre������E[�R�"Y�5��ʜO㦠Ph2���-Ĉ@�OS�8v�b�t̙'O�d��3,9Z���%ϕ�����˰,%��be�Izh�:Г�L���[�O�o�g͕��d�叅���*^�S������@K�r���VS���|�j�a/v"M��tK,��f�vw�?OӞ�*��?����f�/Eh"��i�$<�K�{����>�\	�^w+�a�
=z���u4�|�b�v�Oy�R&����N���ʬ���������������U!���g81���[ka%Ѣ���c����7�p�]y
|S	9��d���]n�H@ēv��b���]�JC�~�&�����N�7{E�R(,�d�p7���T���<f"��IP�6��jԜ=}�ӝ��|�jk��>ЋIj��f�1�/\i�N�)A>F���5��/�7�D��Ἁ�-{�h�>zc�[��dʡ��Qk3�=�ȋ&<��x��gq*��#\� '�2�
���6�Ɖ:�<Ær1oաͬ�9�ɘ�-~���oi�z[�e���2#��ː��$�א��=����i �vğ�09Z�W��'��Fe����6�u����[���w��'[�9n�`ֆFS�����2�Ԇ��	wIo)��'IA�"A"���>{߀y�x��{������ϻ���J���a.����I��!�#!ZB4:�q�b���
U�����l����ϛ��Z����f�N��|��;�y�!�~�^E2i~���[PP��MV^�5'ڗ~	�v����D#�V�@�h�w�9��{�X4�i�k���]\%-��>?Ƒ�e�W�B̘�U�^QM�gDr��S�w�I���!]Ӷ�Tn�Fw=����2�i�(�:�4mV;�nE��+�j�A�!��ҡ��abr�Ƃ�%�� �_�Ղ��WO�k��&����)����^nf\�Y�B�n�h}:�d\b�H+g̥�D�b��0��f`�88���ׇ��.{�R4��ꗈw%!��)�'MA��:VU�J5{qQv�x�[��c-��0*�G-D�m���Wg�S�ibU��<�?�IN�9��1�,ܗ�T0��HZ{��}�b����sCB�jݎ荸i�P�T��lP�>Q�}*#Da�)"�+H���f�_a��Q�R)�k�E'A$O��e\ ե��u'V��� ��(�?`xƢ0�Ls����-�B����|Q'�ډhe�^I��ҹ��.�³�E���0��ey�o� ��¸���Po���R�g�+Ґw��f$Ჹ��z�];Ox�4�e�qb
��E�Q�>����ڐ�����+p�/�s��J�=pnB:8˛LIॺ `�ǈ>�UD�>��o��Ȝ
]�COQ�w`��k�yvi����_{�V�p�6���D��!�H.�2Ҍ5�(Yw<vw�U8g#2�V��"$�A�Z����h�����}�6�cT��$�`��~�_� ���}-�[�����f��e�*��!��p���Y=�0,d��I��(���!�E��O{c��
��'}XI�)M,w�o0]:UV(�z�S���>�Ǡ# �W����db03v��o�$5���%v��R�E��g�[�f�Fu�>k�~���6�*�2)�x�|��<	�u�� �v�|��o蕵>b`���H^u-�Z��)%<�.���������0c�y�+SQV�����B��V-��i�~�!4�d'q
�����'Q�?�_FD�ix,_W]�.�.�.�^��}����U����B�[ُ=�X�,�/��K߮~�ȾN��-�!7�Y���vw" ��վu���#�2�'�T]qeD׸�E�*���Z��b�k}�s{�_+�ޤ ��x����J�����m��ܖ��n�ͬ�$�}�t<��3I�L2�߳�F�9�>�0 q����� c��LZeN���b�JԵ,�S�LF��(���Y���Jf���#�w����UY0ᆠf؇�&�' ��v�ʋ�.|��},VC��=�*�ĝ��
'N�{����A�ٔs/ƈ7ΰRF��p��`���%�m��bp�����ez2��# ġ�C��\���}�#.!|m[�F{"���B�x!f��ݗ�6fx�HǈGG�i���Dz�s���v<�?��f_������hY:�Eň��1��[,�:;�����QZ�P�?u����2� ח����&n�2��Y&�k���������d���>��u(�!;R�L5�`Ȅ�c;�m�|G��_ѫ^4��Z,z���[�}i��5��U��G�Ԟ����jq�ī a��D���-�%�p�8�҂�xhMۄ̢�
$k�$qS�!��� ���Ӟԣa�=<�8@133��B��@�>��&п�e��	Jp� >1��0rcʫ!S��D>�|W2c�-�^9���ޥ��'�7�$5-*�Zi8Un�T���yҸrjn�YӸ@��t���U��*�Y5���c�g2Zn��Y��!�#���$67pE�O��!�?n�I�H;;���$5�M(9j�Ȓ&*��hzo��od8a��\��d6���A���¥-�nw���**��A?��1����i1Ch�,m�F)���ܜ6Of���f|�&V�L�}�=�U����S����J
�Z[q\������>�/��ַP-�,�X��ܗ�zL��/8����^~]��Dl;���j���oYRV�w�֎�tKc���� W8��J�Ns+���Ꝥ)��I׳DP79.$�O)_󟍓q[���[�c���-��������l6<r�BM��r�RL$��PY�6痃���+�k��-�&%*��k-���hg�����#��s��n�-x�4C�n��^�Y��h�/xm+&1&@AL|�[c����cb�O�\+xh�E�n�/6��(��BB*�)�ۮz�z.�=@�\��kK&m�-Li���c���,{}8<�� *��*��&�wTd�d�N�SKT���TCR"�cgވ`��2Hh��xqz3c{���P\h6ȣ�V����\˧�h���� ���~mM[J@����W���%�mՑR�����j��L���Ԡ(Lm�_����vZ�L�`j%;�TT��7�b�*��u �h=�È4������ce�A�^0��t"N�h��߱��-Z_����X��S�8���To�^�^���H���� �*O1�,�I�HPk?���KO)�gTO6�����J����I�����L�t��9��D���|E���ikBM���!�	��M�+f���F�OP���o��#����YQ�ܾ�E�;[���|��\4�s�p��ᚺ�	9~1�������i���	�����1�K�V��/��~���E��m}I(��޵ԛ�l��aa��N;���:���y���=:��: Y���;�[���ĩ_�:S�cuq� n �������)�'����m��#����.�TwF��˱\��=���T1K�����H&�Y?�)���V��[K�P�ɉ���}�����YE�&D�Q%0�x���TרL�x;�ZC Sw�r�|��B������b\�֫�/�B8g���N)Xzk-�LG�ҢPq���ɪCj�E�g��Z�q~$�����
�9L��	��C�4y��ɼ���6F�DIȸ@�t�;�jr?m�������^��Xt�A�Ul0C�!��a����| ���ӡCV��OުNɊ>;��Y��Ĺ\�8����`��#޲��vxR`����&, �Kt�'�\�C6�j�s,&(�.zl}�)�Ehwę�E_nn�jG�of��Ew��<�BJ�t����;˟Iz�Ӎ�{�z'���Y�;��;�,��P��ez.���j�y�(URY)'-��cm�݋��{r���K�iӄYiT��m_u���>�Co�+�a�Q�C���I��6q���C�AyQIɇ����$.�R�;�f�������מ7�x��"���hEfdP�Qؑm��ܼS"�����66{GD���ł#k;��Fx9�!��p �wK����66ofF�ǹ(��e�e_��[�����]����`������R�
�v�Շ�%tz�߭w��&>��i�������ƦΈ+p����ڤJ:4|�ʰlu3*��?[��M�G)q�S/��	�r���g�J���"5�4Ec�)'�!$�Ρ���.^2UNB���BNH�g���L��q�� �E�rmJ�����hR<K����2m�u������`� ����FOݻ�n����O�=($Qc�wV�o[=jc�=��a�z�T�z�4�8�_(`}��~+�E0oJu����L^��s�=���X�E������9�Bm���j�_kjx�ns������M|�t&r���gc>��P���4�s�ؿAo��Ton����>l/����?iZt ��;���L�ǫwf��G:�۔l_w��?�(YƮ�`°��R�ԢQ�#Vk#�͆��wk��6�*�6}.O�-��d�s��{	��m�$X1dihxt.��8X��0�@�i�}��#؞����.�������GX���=?^Naa����"�6�b�Hn��`�_���2	��QR�n�b��ϣ�k�G8ᏽۏ�^7����à�3Y읫�`���/P�"X��lc+��{�h9tQ����[��d�뷣ԧ	�NzB�4�gIH����-�(�Ǣ���L����/�62�3���ꏋY�r�;f�^�6k�d���'���K��[=9k~i�J�;W8�p��{w�� IVV���|��܃h�b�Y,���� �Um#f�\���K���I���E
�(�����i�dx���Gp�9�q�^�����|����U��`$���Zrj�G�;�GNNZ�I5sV�ScftI�����̩���=�S_g�v�L��$!����@�g:��o5���+��]R8F�%a/�S�!!�G;�P"�[�c4i�s�w�L@d?�J�A�E	��/��k���EZ��H1�cѸ}���]!b�xr7_y߳DĂ(�#F�uf��>.�.��O	�V���䎧����:��>����Ix�Q1@Leo*��"x���)���ҡ�^�0��@FHI	�{b�(�����Sy2G?��t ���.��������~\�5=�m싂��嘫a�����AB�E�X߱e�7��J��e���R�Q���JFڊ�;�fz�z������^R1ȹ���w+�;��T�Mf.*.~����i"ٛ��̓���"�q/R4{fWTDC��';3��Ѡ{��Z��L*3���11{�m�z�h $ѻA?΃�$[7�j3�֭���/	�!��ɚ��%(����s.M�����b'y�ϤX	O���]%�Y������=�v��O��_����74��]�s�P���ȩTV�SS��by�a�I:�n�r�X�3������Dh���2#�_��bP�<W��(L����ᦊD�y���ӄ�|�߅����(�)`��4q꥖ʉ����w��a�	���]\��̅��W��Q���K����f��ph$GCC�i��vuw�5���*ȱ��YO�, |�,���|`�+�����1�U�����ޖDT��}��6K�"���1��V��]���{n��;���8�j��]ޜʅG�1gWE�5R몈t���]��=tk3.�K��B����p����7�sT���i7 y:�����617���;ΒT{z`����72�Q�Ď��\�[[�s��p��Z��,D�����W�ίƈB���/�{4���4��R�A�А�a��O�L�v���Ui�*///ZOccg'���G�$Ӱ�E�-:O>�t��5o����+�劅vs� A�.��/�2r4h�B,	ڍQZC�U?�Lй����'|�d6(�51CT�F�9M���"ܯ)_���ۏ�}�4_�qn/�
FCS+]�bx�S��\)TQHMx��j���c;H8gU�@ق�?EU�� ��t�[�<>���P��j�?z��N455�ʷg������˝?�sbM�RE��r�;�a��\��Y(�
vx��#�`�V4��p<V�s挼)A_�/�Q�E�B!��S��K��H��;�ܦ�����5�K)�lN]s���i�
9�;Ə|d��/��}~r��64��i0�y9�TV��$ȫ�ʩ�DW���]�7��a��;;W���@-��[�#�(<�#�&�k�����fҋ���B�$?ŉ�9n���vd��R���L5p�����2Y�z2�LgP��J�mwtNN�pDa�֒6n���G������q._�Z�t�t�^�l����R�m�
�>禶	
����
ٹ����ȪyW�S�'
tT��wU���B֥���v��^�R{���;n�{1p��+�K$
љ�fEN�7��X*�ggs����y9C�!��y�g�&U�hʸ��$yH�U������L��7H��H;d�VQkO�)%H� ˥}�(��q��Sg�n��*��|}}���Q���E�~��a���dk#VФ����XqF��G�yd6l/��������AAx�G��p�ҒI���J(fA�X�y��-�-���Q���G˘���g~l�Ӡ�rQ�+*�=~)ul�H-�gهA8�i�����P��"���đ��o��������_�%�
.�,� �^�&���gfM'���L�ɀ�f��p�̬��d^����bd�{��L�N6�J���0t�Q�'�$�!?D��������6ȋ��!ۼ[�.pn���m�d�}a`��w�,������m�=�;&�&�oC�L�Q/gM�!"�������=������8H���28N����b�oⵆ�?o�g��>3�3�KJ��1A�}}�����e�@��:���Zkb�]h�#��TV��K���?+�a+��Pj��f�N�B�ۚm���'�H~J�HL�1�$���-/��x	ٵ@�Rr�9J�%2LU����l�ts����g�VH��4�]��O�zA�8n�#M���2(�AWBnM�.� T�>���p#��Ņ���vѐ7t��_���}3�J��htE��c{ß��B{�ji��i�r�!�4���~ �Ny�M����&�*���^�\���:{��4���;��pJ��*M��g�#Zd|&��A���3q��)�����>M�@u�*<�+���t&K��2�,%$��p,��l���ƶ�������ZR�tlo���:aB��(|J��=�L;�P\sr���9�ˤ�m��	���qP�s1Q�s���n?eA�S왶Ω��ӹ3���`�o�/��q�W1�R+��)�����_��d�W׏n8jNu��P$MB�U<|m3���'��+	)��i��C��¢_�����]agRӮ���vW(W)9ܓ��p���Q�6�< Oy	�m��C��D�ça�2^���M��W������0b8tؔ=8���h�p�����3�i#�쓁 %��6�{bez��	��8��o7����G�\ �Z�)w����������M��O�f�o
��~d�us�th����UZ�֚�w���3�������(��� ���i�k	�	�ŋY�����E?�ǑWkT�� �_��f_XrWy��-��ť�¥	����]���O�6ӊ�۱FK,0��y�U���+v�o��-0)>4�,5��,�F
E�")���h���|����-�l�����ұu�P��e��#�ņ�6%"8]8��F���ȜF;��H�6�����5aǿ�G=ʓ��t��o&���C{ ��<69}̆�֩���r4�Z�γ�!?��}�&�J���o�˔U�j���n�t5d���;� �,�/��q*�s`��ש�q�(�x�]h�C]�&�fn�.&��kě��	��f~�vc6��gtkːB�>�ٽl��$�������������{f
�	��;g&�T0��vNj"f9�P9@h6����2\h ����Hؖ��E,�lw?�6mm@�Ɩ�*����1뫛(;�*Q�l!<���~��E(����Or'Є�+��ޡ��v���Ҵ���yA��,ڱ�Żq�ab�/�8˅�Yt�,-Sf�8���ȉG�C��un�}ZuWNv�W�+���ԡd`ʹ��PA����,`�c�&\b�����`*���嫉`�҇��E���"����Ei�onL8:l?�@� }�cÄ�t��A�nU� `F�^{�w�Z�ͬHy�� XG2���n����xsq>j�F�c }C�D��V+�gֱ�W^��}�ϫ$��@�Қփ5~�]~��
:�kƑXTk=�D�5�
,|�%g��}Tb�ɥ'$ږ�8�������3�tH�\}������v U��Z50M�#M�v;{�׷��^�.��{$Gլu?�:G�i�_8U�|Θ���W�ՌM~��	8���?Аav�Jf�W�K�$�R���:7��L�镍:��I�.�}�߰:I��>Z��pW���^��	��Mzy�� ���_w�l�r�ƀ�����l,<�����W��T���ޠ���?C�HQ��u����2���f�P׈&����zb�,R���m<��%�R�o)�}$#�@��$Ʊq�F"�F�	�X�����|���:҇�r�k����"���rC(�I������>>) �
��ѣ�>þ��	*"�}��\�p���"�%H��>�|�< �+��~e���3��#��R�5������3Q]mC��<��������ݏI��̛I�@v@7�rK1 ��M���ZI�o�"��W"J�'g���5I�ON��$��{8�"�v�!�����&�e��v�Z���O�����\��e�e ���Y�QW��S�xg��9l�-��!I�4r���D;���}|m$��/��<<�yD����`��Co�@[K#��R�<"�Y�JzN��$2yɘ����?�g -��ta-�e�p�T�9�Cd��x1��\I]s����3��ln������*)Ɉ[!&�V���3�-��s��mǣ�m�sϸR-��$U�xe-��ԑ]=P��b���#����2�JB��0C"I���y�.Ο�{��n,}-f�� Q�ڰ,q�ŗjI�W��م����p�|���|`��?5�3&/��C��%_"x�F���:�Bϩ���N���;���B�r�ۧ�:��'f�Y��P�>��$�.��u�� ��,x������ ��9���4�caL��=w�^F �=���ׅI��W�MK����Y���`�%�Vx%(t�2�{�����'R1n"�
[��|��I|y�W���B�->�g���w���
�II�|�3��� a@=����u��%eX�9=� �u�h���g�r\�d�	�+�f��n@�[} '$b�!;��5g�,>�v`}��Z8I�G��R�� �߂|�V��5���`v2 5fl���b �&��zn��HP�����Ȥ���Sԉ��`0�/��N�Ҫ��?���AJE�g$?35e-�l��:��+fmr� n��P����g�@����ƏD�m�_�y/X}i&�a��:�E)b�y������)�J�d%��t)�ȨY�Ñ��<D� �e����3��/N_���l��t�f@&H`h_}.�����FpL_ݱ�(G�N�������Z�mR)�rhA�#�iةcE�����O��tI��C"B��	 ���e��p�b�c��v�F���Y�Rʅ��9�j5����|�ϡ���⟃�	������@�9���}��N�@��[����>�x$$�ZĻ �{컇���X�id�n� �U���S#���𮰪b;
��^�H!�9�y�n`���K�vq��|=���uzA�B�A�M �"�
I��R-%��)�������g���x������XC��ǽ�9��ګ������%1کEv�E8�8o�/>��(�/��^4[V���ھ<yh(�[]�1��4�^x���Gӄ����ҭ}�9�h�,� ��4��8�?
L�Q	��an4��߫�:oGu9��f����q�gǑz�82��H3�Ip�ZK�'�R�F�N8������>�VC�����k1e*=�kf0џz��YC�zI�����"����ib�����U��j�����I׵���4�`��jtV�M��И��Q|)/�_��]���vJ��\�+\}(���7w.��3��8g�a��q}EF���e}5���������1�mwT�p�d+�����,̓P�i����z&2U��>�ɰ�� �+�oA=��9�r���M��J�{_þ6d9j3�ߖ���85^<s��z�{�7#��*���Pb���!��9��z�&�k��A?���mٹ'�rV��Iy�4�_�[�&7ԅ��~S����zID����s|C����4��'v?���O1ڕ�1�bl�����u^H���8y_n�L�e�B�^��8@��Ta@~VN� ���[�XX���&�� �Z�>�WE�Y���PK���F.��Zz��U����+>zՔ��~��}��X�͈�;I�τ�V�+�v|����6���}ق#U�Q�a
2*o+���� PK   ���X����+  J  /   images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.png�WW0 �]-�+D��DM6DKV�Ѣ����Al"�Z���$z����:��V!z�������g�=3w���=�:Z*T��  ����[��E6ٝ�L]�{K@OUco ��� �����|�`>z>k/{ ����x�Z{�xx9��J=  @Sj�r�o3v́�I�L��S�g@`
�\���EG�T<e!�����DʲϘ��|���E-	:3עt�&^7Cx�-��
H%TH��!�U����������C��ח��(���~�|����>��`����e�~�L����E`"#�n�����bng��0�d�w��f��u���R?	X_�B����������`؂v�r��I���ӑ1��ԙ��*3~��_��:a���skZ8��[;��"���� ���p�HZ�������1�d���g/ǚxx���L�	K��%y&�Zt�Q�� PKI�!����O�Z��k�>)�|yX@8ҳ�́ߖ�N��+a�i��?���m�ޢ�[e�O�M�����"si�n�4{f�g��!l�4eqz� 4W �J��(����3=�ͤ�;[AI=�� �Z�G�'�Ci�55���T�eqo�Z�K��T���/���m�p��&�5��(��sց�ѽ��;�:���v��F3��� 氉2��G�;H��1��"�{I6WY�#�JJJZZo����gKJ]����p�Y�*�`��&���i��&�k}pp���F�oʡ�t ���>�x���n�3c�ºk�����Vq�[˛���ai�ɢ�L�7~@�ĩb5�W����`S�O�=�\"�����j��oq[��Z�ޛ��~z�G��/��G��)����Ci�h�k����i{(z��_�zģҕSD�i�����SO���"҉5\�^QY�u��6W-"RoMaJ�`:��󸼝�@�&�GH(��3wkװH<2�wgv�9���>�M(�Ѱܢ�k	u��WKJN>��`�i�꒬����Bfxn'�R��c`P1o�9��T��E̵��h�ޑ�OZO��F~��nL,"�h��UO�����`�}�p�P$v�"%Ʈ�Y7;�>��B��Q�2��'�З��>Q���ߨ�|��>SU &N	�}�C��<&�uDi�ƴ'�5_��i��H��dƱ\�7�[�i�^�6WŊ6G�M*U����o�c|��3��g��4jf4�퀋�Da���B�h�bs�H��Lu���_b}���p��9�ib�h�Hm���I���� ��w~�:�Ǚ��(�Z���iaa��-%�X�0n���4�S�P+ҙ=ߊ����D��BmvI�Mm>���}K��A�U���q���LyKHk&��MjB��}���A�f�)���D}�ü����{����h���xܞJ�tW�&P=�a�kw�m_,#����rׇ�߶<J��V�vg���^���ҵO4 ����l�IGB��L��PS��ڽ�����	�;m�y�}a�.��%\o�jͧ�g�# lF�<���s\RCj�ch.�5O</[ߖR�̔��{o�Zwu��H�UV�E���_�#>��N����1�+��Ġ�E٫�ͺ���vub��Vt���9c�M�j]�򏻏aj�(p$v&�99�r�ئ(��J��Y&躙l��u-�1�}x9��x�=Y��絗�<D���T͢Mxf6���Ȉo�����{�W�������fF��Oʁ�����w�7���C�f�<�{a��ḡ|̴n����*��V̶Q�$��e���YWc8���dO΍��$V� =�z�z��!�Nj��8�H|������~@�����;/4��ʽ}�Btnb��D��WsV�_዁�tPY"ۃ�t�����P��~/�9žcT��bQ�F���n�}kM�F=��(&�����<�{�W���i�1Ӣ3F\QJ�"�i3���%��1�ixjF��aƓ��r�*:H�s�Q�"�@�g�����������$-x��d�۴�D,hO$LDRS{�T����ib�7�G6CK/X���7�ɣ� �)��֚��tWDE��+�9��R�dV\�Ѽ����E���X�;+�[���P�a�Ze�J-s3�~v#sA�;~�sDh	.l�//��ܦ�:�S���Ż��|������ᬹ��FO�����h1 W�f�V��e%����\+C�p��T�8�wʄ1���l�5k�a6�|z��j��������2�zX��:�ϳ9	���P�������@�UlA��0Ԥ����\[j�4�r4�j:UOz����'y)c5�����;�u.S�����t�i��p�*y�0ؾT;bg2015A?�Wj�l��ۢ�$1ye��K�����E�^-����T0���8��� ��p��a
�`h*�Nj`���S�^N���dB�@#�*N�CK����9���R���૕V��v@cy�;�K��z/:�,Xi6S|��궣���M��v]�� &)��\�4���9h����_T����,��u��=�n2�O�R$گ�[?&̽�W���'����>�޸��R��q�ݐsW�t�)���9RqP�`��]�
� }5
B����g	k��g��wf�Hf�1bt��}����8��c�N,���.��)��֩LS ���5���梓EjP�r
|-�������q����F�(���5,�y@� g���Z WMP�;�,8#�]$.%'g�^��!��.�x-z�\��������NQ�{�zAz���Qr�����-wT�1�,T��r��5:}�R��`Ha�ځ_��K��������`��s7}��3���ڑ_�129kzV�0��� ;�#+w7�p�i���L������ xT{�^W(qm���_N@xGY׿�<�F�^�FNz079[WE�D����i5��n����a�Į<�={�ܕ���V�i���ܬ�K��$�GȰ��ץ8IU5�D:9��W�Ռ�,!���%l{)�8Do�P�H�~5(�\@��S�mmu�e�m�ڥs��>+��ڃ	:=s�Cl���Q�X�f	Ǒ�V��a�<Z�5#u&r8▴ ���c����~��?�j����Q�EB���C��C:��h��a��L�І������l�z,.���'1yiV���F?��K��.ϱ����"�lC�&A�{>�v݂���`Ԏ��:���<��Pj(_�q�e�E}��*Sy�ţ��)�E��k�����N>�a��Ȼ�U�Mċys|���_�֕�d�.#pѫ��4d1�&@�h�[�Q�����仚b.��W����M��R�k9�FY=�t�fn<O%����\j�l���t�r+�����Ñ��T�(E�@D�����3jbT��hy��b��A�`j	�\)�v0�	Ăl�r]�_��_�%K��*����d�PS���ſɅ�.��{ӕ�#�X���b�\6��K�g��,id�dQ7�o�|#�p���JN��w��
F�$L���2-x�s��`�
�,"#���ށ��1'Э��x>���
#����-�|a�M��^Zօ�Q����q��>��Ւ����v�Ur ,��[���t���(dN��z*�Vvq��}zR���j�fC�;<he>��4�d�R��f�Jso���|���_����|	.���۷�R1?����#�<=���	�of�d���{�-����k}2`Q�5�����/���q���w���t�B��a�˳� N��%y�{�es!}̰B�crY�	5C���ņ-5+z �!�K��U��9i��hE��������$M:a��Y�UmW���JU������R���)�\�Z�~[O��-#���b���T��\p�������O���h�_�fR��L�����WNs��B����z���{Xc"]���oMe�X-��sī�M�`��E������[���Y�T��0�:������ϟ?�=�
^p�>f��ݚ�4v1>�^���f��"ȴ0��^�f���J�j�M�ZŐS_B�M�/�������c;��[�sCT��#�܆���b���?PK   ���X��_8
  3
  /   images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.png3
���PNG

   IHDR   d   .   �!�^   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  	�IDATx��\klW>3���?�vR�ql7M���aBih 	�F4��hS���H�

�U���u� ��[�(!IqS�R�j�4&�;i�:[�w׻���|wv���cg/�u�I��uw����{�w�4`H�b濙%�k
�ٟn�N�W�éR6���KCCC�v�����$I��$���|�aM�<p�@ʿ�Al@2vPq�	�L��᠎�jii���2ڲe�,��,��=�}��7�~�o�.>��~��Cs���\AY�)�1::J�XL�c+���b����0E�Q\n`6�?a�Z̜	[w�\��4�
�"���(JB��|>��}\��y���y�j�̝�h��t1 ��������X��rrr�6�������i��̏2�j����ee��UUUTQQ!���A�Xyyy
�(>ȧIp�bA� Q�������w�gQdvk޴��;�oN�G9��9c�ڲ��1��Ջ�x��^E�2�� vݫ���vH*�Y3J#
��Sv�y�F���|
!HT��By,�|�{�1J��i�D��O1ױuT�y|բ��j^ՈcwH�V���RJ��@.i'Iי ��L*H��ͤ�wyh��3�PN�������v�j�**b$}�O���#� 0ہ�����TZZJK�.�lc� �������137~��	�Ht٫ju��+�Q%���3�|��a[Hz�$������Vjnna�֭[iѢE��OD�@�c������������Gn�;�>�Z*�B�QP���u��r¯�����cتjz�p���OИ]�/3_3��_�����0��3�K7!ǝ�xvb4O`η�3��"��V|ְ�y1Q9n�O4M�.]ҷ
�"�"��0�M7� 1�a�$������h�8.o6j�0m�{�<y7P���'�lo&c��Y3���#�1����9,b �:Dzd���drG6� ��O7j��41NG"#�L��Z�4>:zs���H�̤�1�!e�?�>�|��b\�)��{|k����8v�#
`�:��ac.$a1�1Ě����2_$}�`��[�P
b��LwWf!�a	��T.m&� c�
��b��(�1TU�'��nJ#YɎ@" ����I�������@�������7m!�8�m�9XFB�|�]�{�r|����5 �h���T��)�!_���b!L��_YYI۶m�ˮ�>����0�}�k���N�ec>�l�J��'_M�ҫV]UN��������~����w���"d����.^�H�+J� 4���Lit��g�-[�M�����A!�����g�v�|����vwM�I�i��)~�9��(+$g]�k&��+W��,)�U!Z� �"����療��D6`%��� 񋵩��O~�܉?z��G���X ��$)\��˺�|�k �������^��h�����C�O0	h3�w�*w�o�N��p�7�Ap��W>L���p��OJ͗Y_t�|����Q޾ig��o�7=!����?�)z ���ڵ�x �or�Oix��a���YN'k�厰�dG؋��\�ѣGi͚5�v�Zۑ�b	�+ H�����-̳�=��)�03qc�AQT�V�Y# Az{{EZ�������S���&-A���I�:YǬa��|��i��	igS�l�1�Ng��|�t�YA,�Ę���Ux�՜G�W����kMY{� v��g?G��g��lG�$��q��MI&K����l�anX�g\%�*c>�\�<��,�F�)D9����R/��]���q�6� �q���"�W��3_���K��9tn��w�F����6�m�K�u-����`��XS�JЩ���1B�G��������n%w���HԈ����{TRT�R��DR�����yqu�0�G�%^�1k�9���+�]��z��8�̿zK,�~�oJ�EXz_گ���JJ�"�d��@�ŋu�m��wۘv�iqa }|q>�t�q?q��v?�_^�����>0Ԑb���Ⳑ�]�z5����e%Is QN2�3�ļ/Fr�S�_�i YEx�~���2��,c�,� �t�b�!�!������"�z��5Q"&Ǥ��b������ҵ@΀�,��&����s�GI�X�e�(��܈��+A��X�`d���&�dd�/�L{�rB��bx����DVbĳ�R��Ф��7���Q�$eOrр񢧵1,���/��%%%�����l�̉ �P��������K�:���6���Z@�c��.
��=Â��g���O/Y��������]�Q�E�\��46�]̇������6k0'Q�}
�Y�v�+W>��Y�h�U��7���\��� ^��z�ϝ:uj!��9s&�����d�?�`]�ḣ��k��(�ǌ�Qbd����-�Ik�S�l�C��%�KX���Й��%vO�g<���شc�aM�a�}�=�
�7    IEND�B`�PK   ���X	�\  \  /   images/898ac7d1-13d0-4a1b-8b5c-ab7066f4327a.png�W�W��%����K`鮥;%����n��I�EV� !݋�t�>��;�̝{��qft�U𰩱  ���"��:��&�ߔ���'X^���  ���q1��w��S2���t���y�s�p��z����T�|M ��)���YfO�����~qv��ّ��v�C�m��� 91��3�,.���3��2м�P%sVOV����$�\09�U,��Ka�����fv�6{{l����c}uu�ڻ����\"�4����h�v�Y�!^����!7�)�Nʑ��[��������y�B�{rrr/[��q�$�|g�Q\P\�_��m����?���Z�|�}�X__�-��pM���������O{uNF����0M8�W-�Դ��۱�茀��4�7�/c���'ˎ�{ƀ������ka��r-�v����}|/}||4�y}>~�w�R1)d�-�uYvW��������kkkW�O��V.nn�� ��|'��I����K$A~���:���0/�j�ڍ>�^�,��ۛ���x��krΖ[�2��������I����}b�t�#���3jL�Tp�f���%�M��&g>���h����Ŝ#)}V�c}pr`�A�W�rm('���� � ���0���7, ZB��{����p_�u~�>55��ŗ�L7u��aMH����euU�򢻋�@q19n�ViFq�{$'��Q2��SGv�< ���Z3?d(9_�S���'���Jߧ�kc���h���dNF��1�;U{�K�����B�~�o��JL��S�d���b��*��+f`uy��[!s^���w����%]�sCã�~�����������x� �r�fr+�T�^����>uMֵ�컁1t���!��Y*��%p�fWD�����Auu�]��E�R999�e���R���M뭡��'�i�=N�#U�LԾ��<�ۯ���g~��d,x�>�-�&Inv]_���]����*V �|�������B��.{��,s5��D���#��Y�]��f�h,�2�@������?@=Y-���犸��{ǦvFϵ{�����eI��<�T�ۮ�?�=����#D@c]�!��Wg�>6���g�T��Tnƻ;� x��ú�(���F�����.Y����֞N�;=��U�v#�Q�EA��� ���o����T�����<�]Ц���P�U�X殎1��ٽ���ş��z��ɿ�eN�]�jGs���\{{�0W�5(���f��,4��S*��A� sIh��Nw2�J�l�ਜ਼��X�2h��3x��%Ǩ�j�L����	!Y�@�G�s��*�l���#�ie�	IM�f�� �����W��D�����<;a�+~"�
z��;B�t�U�ť�&֗ff�1ɭ�}q��2JZ����vj�6q�^ c�Ì�M���(�0E�⇥�<���-��~ �*�塈(-�?���Ć��$??���q�yr!Y��:�	�7�M��m��;e |F]Z0�u��Ӿj\pW()I�+)�F�8epr/a'?�޳����]_А��Y�5�����ff��Eig������G��i�	��7?���y���yVq�]�x����
��1�fs�(�/�s��l�R:-���^(��6?�s���N?���eu�-�&�i�czkH��Q]��"uj�Fz�0��a��5�f�H�EK���c/I{k`��pG��ߥ=n��[����ڥ.w�p�a�a*h4�Vb%F�J�觍��vgc����<n�����a��eG����U���A�5��֊	w)��~��+����i�f��uaΚ�¯��k����[ ��陙�.`ra�AlqC�h����6�S��'i���nSo�'�$���ٹ����WKF~�!��%�0d\��Em�O]䃍��+��qLi�\���k>
;|P��&�Q6P40L:G����J7>0�e+��f�Ԡ���,��{*�$��Q��$h��#��~�i��*	:�R=�0O�!�������d�!8�۠( 4����U��-�l*�L�� ����\���ch�*���bh�J؆*�m K�1��JM;���s��¢k=�{�5���l^6�&cW4|Y}}wl��j�i{�y������Q�S
�	�Jk����rl(@�%ݴ'm�ڕm~�����=�tLV��%0#)��{C��@Z3��h`��[�0$/x�t ��g�?�H�!�B�tV�+61��BG�nna�R���o�^2�J����+�Oic6|������$��,�8`��~K��	K������儃��{(������v�>�)�����'�ςE�\���udJ�HG����5�ؑ\J�M���M����D[���#y���� طt.����Z������C�+[�H�����nK!IG~\���@�#.f[��=�-�#�=	�k�T����B-�m�7��p�������'��9BL�[Xvل��Ԥ0��L�;,K��Rd�n��5���,�J2^�A�+*RR�����g���U�)��ݗU4�����s�c������Fۦ`e�m6vX�t����V��X7��������F�M���1��7?tK�z+~>�\�鑵z���.���il0Ͷ��z�����o�j���W�)���d6p�n��X�����5D���'�((���W�_��r�wu�5��b��ߏ�7{4����۔iA2�x	O��o�ͩr�Alȅ��o��)�?�P���/J��(��)>�-��qQ֒7�������q��a$��7�N#&msܪ��/pѱ3���H굪F�H%n�58��G̮��*�'B�87�����%n�p!=ExC���'�'�F�+�,�2���(w�Q���Y�� Y�XO�Y;�2�����dI/#|�%��z�0%%��=J������8��]�@y�? gnd�ns��O���kI�dv�E���E�/%����@���q�L}@N?:D���,lJ�#˩��fh7zC���[��K�1Æ�5��Y��5�UEd��{V �8�f͙��:P�h9_���%\�}����7�E�P�E���E��1D;I�8}��rO�C��\�&�Z������8{3ͭ�M&ވ
 p�����4�BtuP'^
��/�Q���[�$���%��U7��Ĕ����v�����Z���*�\�W�U���gj���=}���D�hR#��E0��fi�ۑ��>5eY���3viܵ�e�����hA�v\z��7���r؇�ҭM�iPP6ֳ}��=����u����!x/�E�`�%��c�<���,G��
7Ŵl3���}S�A�:1��	�p�����_�ð5=߉|Xj�W-G4�Ҧ4�����[�8���UP@����m}M*�Q�CQ�{�nK+hb�M��զ�Z{m���JM�W���1���7����h��PO��)�y�~�6�{�$U��F 3��U_���h �=�������l_G�R*�MF)'<���H�~V��BI��vp�66.�+up�nf�p�y��ˬ�������%��#Ҿ��� *b?0r�p )�ʮ_FCg�^�u�NkRa�lI5�x@�	Ub?)�Y�����𷌌z�|�<04�'�m�r%h?�c�;�_O��Q��I�F��bW��9`&aL�8�S�I)�P��M�~3���Kx����ދ���2���qc��)v���4Z�p�o��I��	�jk���4��V����V6��2@:\WD�5F%�D��o��پM��g�\�!��@�����[�Qxa��F]����/���mA�zl tG[r,?ɳ��h|f�C�f�xgW���tg���	Q�!� ����<�2���
��S�����uʫ�H�1c ��$7ے�]9iJ%��K��x|H��?�u�R��䥏�~�ꄍ������p..�Y�ܬ�ܨpS{�!N����� ^g5K��;U�|0�.~\�p��Y-8/�ة�{^|�1��жٟ�Z:k�2rc���yrS���\�M�A�ǭu��w{ۗ�)���濆���w��Xw�/��}��6�'�Z
��b�!�|��լ8#��;�o7���i��I[�P}����Ę�-���;ɵ��,�E.r���aUț��j���}9$���LZ��N�����Sw�웩N^7+Q�ZrDoo�n&���.G1`��8C�
�v�Rl~Yk���J?:>F JM=߹5���%��'ב�pB�U����V��Q���&3��]M}��L�؁����Ц@q%���v���ߵ�y$Ϥ w� ��?��unin��}�[C�y���a	t³�{�}�^���T�U74L-��9�U#��!`ƕ4:� fPpF����v�N��z$9�;q9���cO����{�m?Z۬.j���Fw�*�6��k ��A�R  ��N�2Ͱmz�����B�?7&&��g�Q7��p�%Q�p��*��۹M�[.ԉ�xKK�s�4����e��".�1* �0A�Yc2�PH(i6D�w�`bQ eZ�:�tb�y9%<�	, �b�����C��+�a���&ղ����;[K�������`����E	�sy֝�w��E��W���������̃VެGG�S��tך��X�����،�����)�U�<��x���~�ݹ�l��{Sj�w�)�ƺ�a���k������y`eQ΁r^��;J��r�2m�慗B�OQ9%$�&Yj���C��̪0�[�E�^l�k��Y���/'�O@mILdw��h�7�܉2���c��_q�������1c����~��#nY�JB��g&jfE�rP+�" bzC�Øp��x]�U��� �I�����gN�@X�5`/9�䊌,�&��>�<p��s�ǆ���zu�k@���9N�v�o��=�	��y�Z�k�.�>Q���+	�R��igF�̚��T�Ǟ	����<D��7w���vUk��ٔ����*�'��'L�.��-�� q[PV���eOǻ�W�q˒0P������sۢ�V�SY�n"�T�N4@�y�M�ܟi��{f�=E�}|��_��#��2����W/4oT���=B�`H�֙�ɚ��JS:Ed�!e�%`��n���q�v\.��p�p��]�l�(��"�J\𘵾V�v�m��g�B5>�w�'�%� ^p
q�nބx��+��>�f������k�Wj��|��j���o��_�ʈ{K`"��vZ�,�[����=*w��Y�R������i���
��[˵��ж����,�"8�s/�(a���M��;�?Zr7(l��U� � 5<��N5�?�Zxn���~Rx�$}I,�OYQ(���8�-�z^��-$�W������0cg���Z�	ȋ�)��R�dA=͸���z������Y�\�+zl���y��8Ϻ�q�=�����6:8m�R��N���`-�J|�����,��!V#>N��Oq�g_�"t�uU���hX7o�m�i�Rr,L��z�->�#8ÀU�#�	6�s���Q69��&��w~�4�~���VC���� "�����y\U��j(�S�����Σ�Z�X�k�O	�!�$�~Q��X5�fѐ���,�4�#u]�1N�.8F=�Пux���|���(��:'�/C��[<�AVĐ!�j����˧��1���:�
�]�}1��L9�?eۼ2K����l�vr:��{��_�3I�p��P���fۼ	O����(a����w��r������̒I|=�����|K���'wJ1OU�#�AT?�^
q.b���\�kr���͸洘�%�Ct3˨��A�|ؕ��`�� �~�Τ$�-�'[
iXS���J;c�wso�H�=�
�w�HKP�~�^:=�!���B��3'�z��G����Oʑ=<!?]`;
�6�������H�&��5U��,/���P�}��մڢ
3V���\[@�e	O��i̝�KBm]�V9�}22�)�u1z��I���B66)X&�ր��1n ���Ph�ĉ��ۘ���BG�AAa��S}}ɯ�*��I��z���C�;i�F�DV�O�	�GV6F�2<��v�����'�/qK�E(�Wኬ��b>��Jbd<���T<�VJJJis]]p�R���SM����3�rW�����BF���7��!�����x����!w@=l̺�㮌c��*3��ڂ�L�/��"U`�*_�!��?��^�S?�z���I�^E��[�ןb��R�G#��ݎ�]���z@�������]ϣ[Cگ,��j=���j����4ݗ=��ڱ��Tu�:$sy�ab���0d��1�L ����G����5�>9�iزiK�VFQ�f���u��?FSS���X^s��Ja:���?QY�����]ǁ�%��[����n�t���>cd�n���5��e�#n�{~co׼�X�LJ���%��2���W�`�ee*���K0Ȭ��RX}	y�q��/����(���L.,~�{�r�*�Ţh�H@n=w�-�˄M�8�sũ
�Z�1����sqw��5?�mVYuz>��7P\�?5�*l���R���"�<=�j�"���3��ՙ����-$ ����I�7n���b���1g$���i�����9���L/��q�#������&�FFJz3�U(SR�S��y�.��@*�'Q1���X]�./��f*�����'��$::��Q}kY�u!>K��~�K��z6x��0晀k�˻:ݴ�+#x+A�`w7�s�dm��q/ɵ����\�ig �ִZ�$���H)���Hd�g��u��#�.����[S"��u:�
8��k5Б�~�(4�}��iM#�����32y5r�`K���\c���׍���g,�d���qJ(�HDKR�Wuk�WY�
�ym�fg�ؒǽ2SI)W����qȮԒ����+�ϡ�36ZB�!B��V�	�(�dϓ�S�,�g�����g�Ih�Hx��Ȟ��|�b��.8x������+\b��O�	������_�K9f�Ð��n��T-�w�s�Ǻ�奯O�F�e3^�����"X���/)7�z
l�50v^���f� �T��剡��O�Z�'�jJڊM�6Q�PK   ���X�Ƚ׌  �  /   images/9185dcb2-65ea-4de0-8d42-42cedb1b5634.png�x��PNG

   IHDR   d   -   X���   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  IDATx��\�o��ݙ�����uڗ��!Q�Bp�D"��h(U�$B�F_���?�C�JM�!-�А�J�(�U(I��E�|�^$k�w��u{�ݝ���?���gM|}?~3���眹3'֎_�A`$�M!p�8	Q����~��Ql18���gv`��ű�K�Vr���x�p�z�3���rW�y�4�0Ɲ��t��=�r�Ҙ�xq�!4q]&��:׸:/s����Թn�?V̕%�p���:�+3xg�X�@?��Ⱥ�qO�W�t�G�����X�ѳo���Ij��;m�I�Ae�ŰĠaä���	.���'�eV�	C	��h�*��2�z�=.�q�k��I�%WZ�A�KD����rB����'H)��8�{?J����>�9���v�4�'���~��.��7�'`��9F+ o	�'�!p��/e��!i{?�CP����Ij�Ҹ<즺aj;C}��Ǘsݥ��N\₱�ߧ�$ސK�\��G��	y��s���׸��s��%\�I��,� ^�cg���CT���;s���/��e����2f�f�}x;����Q���r�����2	��b�\͘�#���-��pb�w��u6�S��;92���&�}�5L|�,�a��ʚ�K��D1p�eM�H��ugDq�ߣ�[5.W�z�D
!����	q��MB\s%��Zs9ߦ{�/�$��b	ӓ9����M%wk|ao��3�=�)㭱�I��4Me����K�_�%?�q�<��5'��-����Ү_���W��:�of?�˸S@�w�ۻ��~Ϋ�1\��K�
�^=e4��"������W]�r�\�ո�k��書��հÛ�����$����ǰS6�}�������>��ذ�)���Ty�"��])����ZMtXT^��s�V>�q�<C%C�u�2�~󘫕���M5�;s���R^����D����}�s_!�.I��VH����k!�){a���2��0ڔ[���̵��`@��XxL�zp�f�S�7B��"s���q�<σ���ҿ�P��J��h��Ȝ���g.����U�^}Qx��t:��C�Z%�d)�jдЛ�s�1�J!�H F����R�����Ӓ뺈q��U!�M�#���c��"(�Bt��]R*��V }�����H'��t��Q!���xUH~&a�����!١;غ5 CG�4�O4䏱z��אi4)D�Ζ)�L�8:$�U�vQ������:�Gx��x�.��~���n#���q�EA/W�W�H��s��������/�]]T<���}t��.��j�G�E��WX�_�|BE�
���Y�0��/-S���F�]̓����@�1����n���~k��j�ل�C�ޠهđ��CW�c�+��+���\�B��T����8���u<6:.��aYC[q��Z]C�r��X	�z�Z�Z!�Fcr=�/��Ut���q�@�\Ѱ���\�d�\���r�r>jp������!�=w��B��B����`t{c��	��겻�GA��lZ��v}�m��_�Z��v�qb����/�^�B(JKO���'a��iw4���������~zHي+ڮ���E�S>��W󉞻�S*;e�d��vr�-�+�hVXG���f䫊u�S�#�J��Uj�pc��mw|}���l� i�!�x_~=����oܺ*�5��S������q�8N��\����MW;t}c844��'G5���!����}yB����a9F{(?"�_�$9�c�3TC!���
)|�B�O����ؗ��0�W&�RxT�R����s%v�iѥ)��	^�U��=+���0-zJ(���/����R	o|�6��}� �3n�����=zw�G�X�ξ���z0;���<w����4^y� Ο��R�¬����i�C�8��y,U�0��UI�c��W�1��u�Q��\�����p�{`�OO�0Br��V�u�0���\�=�r�9=�Va2^��ͅ	!�sZ4+���w�n������ة�jep��!b�~?�7�՟�{PiѤ ��?�(�*��    IEND�B`�PK   ���X$7h�!  �!  /   images/c6364832-c854-438f-b38b-75bf2a0cd33f.png�!މPNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK   ���X~��a� ٮ /   images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.png\\\S�� Áh���P%�lٲ�LX��,��
BX�Q���%�A@�� �0Leʎ�gb!��b�����p�=��y�sB��#=�=�{ /��E���-��|��@�W�]~�a�<����7x��粅"������	��Q�K��&�����N
%�����p��I���%e^S����iP��`ȓ��P�ej�l�{�y�o�!O!rݢY��بߚ愳����}���r�Wk괡XY?�q�?�üh���!͵�/V��xt�e~fc��	�O��D�:���s��;%!�E.�o���˘��P\hV��rɘ �;����TS��{k����EA�n�Z��2���|��k$8V�p�N���$&��������Q�9�HO�	��T�{���M�*��o��f���̑��M�<�!�f(nQ����P/ h�fvh̜�,`�*�Kp��e�Wc=W*&���s#�pSx���]jr������Y�]`7�핮��jʿ#˰?!!�\Y0jn��D� ���Ȳ���h��87Mr�q|h㡴@~�K���g
�	��Xy6\���J��ځ�ӏ�u#H�u!�}��K�����%%%v�ou�V'���'���$�
����vv:o��Dz����p��r��gD�*������Tc����u&�17Jw-16������p%�8Ec��Nl�B�{Eُ��^�LG4� �s3�Y&Gބ0�F�٨����?l�HIƾ�䦚 Y��q
؜$ȁ�,S���fDz|�e,�q��傆��Vn����@>$2�r$t-�Q����a��o!KʐĦ���H9�mb�����m�Ž�u_���is��=ۚ����1�r�|ϐ�B-a9~X
j�MD��+	��#ҍ�֘	��1//�����")�	p[�e�5���(ۯ�N3�� d�)T�����ɂ:�x�f�h/G���%�����	L�e���fx{���}~~~��J�1Ε6/c�&�
?LDD�˓��3�{����g?�eB���Qsn>��>�2�+Ȯ�\\�1%^�+���q��>�n���R6��]�]z�}B�u\����uv�Y��H/$�W3�
&d��Z��v���#����ї����k̉�����ڱGw4ʂ��W/��� Ɖ��OP��m�*�E"7f�TU�����a�@���+���=�o�a5sTL̖=),�Ek�k�:V�[o�_�#� �zbўׯ�o��Z�Wud��x��CU/��Z��,L�s�ŉ�kY�����"NN�9�s?���ma�����i�-g�1����H$_g���d#0[��n�����S�Y� ���>snBj���ݗqt2�0�׏�΁J�����7Z�|�2��_���R�t��� p��Sй9;��q`;6����@��VhS���[�0��o��V�e�_|B���l\�Qq���So��D�����[�m�~��B��D,|x*.F�Ƭ_�8��J$�Asp�y�f
<�]U6��Ka����n�����#	,�~��=w'H�g`��w�z�<s��@���Y�Y��F���#����e^w ^*����&���'�
o��$5�8����j�����	^�,-�%z�h���K`�kʋ��Z��**����J`�W	����5��#��i���h!����6Q�#l\Q�¾��%I�>}����t�=y�y��~pyĒ;�H�Xc�u���޽{ͨv! C'����|SE��u@��;�u6.^��~pG��
� �ژ�m�@[�:�������EEE����G������b?�*���������6��7)%�iv֣j�kP~�Ӑ.�Ă���:�tD�B|{B�B��Ǭ�A���*�m^Y	R���_
�~�VP@���1���(g���l����ˤ�E��m6����@��:9߹���п�YL	�i:��fdZ�c�Z-Eջuee�KY]���mUCEUUF�VT����206.���J޲DvM�d�|�v�3l/��i���9����ϴ��Yy���3�;ǲ���9����vnHa��zC���d�?�{w~��|2����r��,D@���ͫ�P�[�kᅠ�,1z3��@Sd��o�<��Z�x��Ey��(韤�����H@n��̮��0���k���TM����PSc���q�h��m(�Y�
-!��a�؄c�o{�����;Ϫ lv�R�
�eXR9N��6��c�ݽ�j�y묬,�/����bF�a���؉����7��Bl=h����>�n��P�J$�\@���P�y�m����_g.$%'7JTc�e�NLִ����������=�g�'?6�L��U��N��=��g�j4B�- %�O��@%���7U+D���oM�"\�"$�p�� {��+#1���G��P������G�8�f^U� �!߆P��ɲ=�Lb�ض�>6ʎ5��-�m��X�7�E��EvQ�K����(�����- E��ռ�*���к�01>�s��� ')���.Nb��̔�98�p@��b���w�X ~*lD���w��-����B�@�=v,Wc��=�M//Y�o�+����R�U���^_�&�}0sD6�h�I#ql]E"k�뾤�bS�4�]��IU�l[�I��^�7���z�5M�뱂��@��l�wTh���8�4i=8�j|�ߛ�8I��
��$�
�}�{<ڄ�o7�C�+S�$�qU#�3�FFF�����r��ၞ�Wz1��c�N�M�cQ����}�".��O����*m��A_��o
GϚ х�ie	+��dH����Q�kE=$��m�2�0E��趖�`;���8�31J���̧(3�ۅ���w���J/�:��K�\��"��PGe�m��=,����Cj!��W�cVXU��L||*�'d@��������Z�2_9�^uj�B�.+��!1���RݡY����)�&)>�B�פ��HkU��k`"�c�/�oS"���ʦ��6C,��x`����vb^�p�`�Q�Ǔ\lsDY�x�,P/}��r�-i���Y���5dx�w8���t���6�#�q�n:��������f�de��=�����Ĥ6)3=A��\&�x(�EE�f�z�����FWG�l�2�����0�㥒���E�i�^��QV^*S� B��Uqк����P�zK�'T��I|���	Tb�&��S����<��51��W�H$5��(�>nV��*
x�Nh��@�/DDD�$n�'5!����<y`3����l/`���O-P�>��-4�һ�e�U|�\�
�-<idd���v�Çw�����<��[��Fj�f��������L��Ӭ�\�:a���E��)hȵ��Չa���J-���`�[0,�)����
\[��&�,5U�����JT��;6�6	)���/�^�� ��gz�s������]��`w
Q���J�����>abA��V���rkʳg�)��:�����wL�^����6�� TT��B�b���9p٫u��ۭl���2��C�uX���_#	���ڴ������c0�N�����{�����J�H�(�aԏ�Ƥ[����ϧ� T���n.I������;�F)rh���bi�
�Cܝ�޽ks��qF�G��W��9�o/�W�Rm�F������'�m�(&�M�h��z�4�0��z�n�<A���(o���]��4����a�<�$@�V ��om���Ź����+X��H��ޜ��P���~P#ʸe 7�v/��k�4Tj��gߝ���8D>a.�`aiY58ƌoP��UO3���f�ח��/K�j�n*�{�� �@Bv��πn����w-9�E�mL����S��0��/.���WN��_��H�&X����Hnz:�:;CσT�����ׯ_����ۧ��V����K�G�۹��K��>-���f懧o�v5�h>@��'3�a������f�ֽk�mv�G<�S>s�С�xĪ���J�Z��M��k𙅅�)����6 s���1K�^��@�z��ʵ�*�P������"7�rͽ����S���q͹!5`*�/Nu�n8�+��4`�0>֤?<������[+�/�?^\{�9�F㾲�N�R�������d��Ҳq}-kS���sֶ&t�ߟ���N rMJM��Q(:]|��}J[��r+�G�	]�E��]\�JlJ����5��2���o+���T���|�j�R��F�Q����v�\x���%cn&�'l�nP܉��X��М`��C�����Mq�ي�@hz�`�KЪ�,��Y�{�III�2̭mlFD����g�*,�3�=3�X�ؠ��i�y��0I�����P�0�v��qUI��.zn�p�f ��a㬉h59�f�~�P�`(�	��D������,J�`Y��G���T �a���c�7NY�{��S�;�e����3lgL� �s{N�>����$�5NN�Y�%@X��E��A�L�`��``` }����?}��xWt,		��8�
`;��	,���NM��W�^��	�`��v_[��xK���Z�
Y����W���eƒ�@�;���+X�\��XfyTX���C�꼩�o�gwk��oS��I�/����ơo��Y��Ü"1�<�"Q���_�|^�����TSZf{K���kEӌ�'�2j-o����������n�9��ھ��(M=�%#T�c��
V��%�!0ܲ�ܜn�*�ӛ�|�`Y��� ֓�Y�?��-S	�t�&r�K11R�Q֊ ���V )P�L`�����tn�O�֏�#K��bmY���Wy��`�:��#֌mpE銰ʗ��1�!'+�i���>��Y��tT���@�`"k[��%�2����0�nG��L \X�x5���u��4�3 V��`h[�V�L�ri�{K�Q~�E�1\�7�LykMU��+ �Z0��tʷg\Ē�ءj}	DrL�45SY��]�i������B�,B5x�s|�����5�!	����jz���?���m������	�X���2�JF�Vh��>���`靵�_X]��f%��}vu��o $�}���6��r5q /,�Fy��N���<a�
���xS�K��4  \�C5��r��/7|f�}�U���ɞz���Z���Y[�]_�ե ��߿GIlMȌ�p@〩L_�0��r��џ<M��}ZV��5RO8�t��.�@�w&E�_X�Z�T�,,\[����@�W���M@稠`Uy���7����h�b�S?��G��B9����~�e7��@�)���������]s��a��Z�u�z�$�{��$3$�����COh����ۦ���i#p���&J�!�;�\���f?i������E��M�gj��7�OH��d�rйN �`?�Z��x�%)[;�n`����O7=����޵��Ngg��_6���~�rq��'&ZӚ@S�N~|�8&�v�'��c]��K�W��1��4r�	�\<7��Z���߯�>��X���IFݯ�mۿ�l�.k;���!	� }	��3�zr�{��]�"p���2X]3����5�N���K��-��ɩ�[k`�Nͬ2�PXo*���r�y��P��M�A�Sk@��=d���*�D.��'{�Hl,��A�� *��.=�zs0̑�e�oQaO2@���U��o�,� N�wG��Q�'V_{s̰�Ƀ���6�⥒ң��������6�@ث����#|pI�e�(��	8k_�g���C-tտ6<�'�W_�p�ڡ���YAM��&�jSب��}�_J烜��X���l���S�n�%� bSk�P�1ߟ �he��X����<��7? ա�8��J���X����k��<^㲭i"��۱���S�A�M�T#rrr�D ?ы�\g~�(QQ�fV��O%���,6腟g��K`��<���s90���4X?�B=����/,���~�2y�a�[�� /Wל���!UY6y~ڴ���4$�J������u�g���W�}�8Q;^rݹ���%ǟoO�z���U�}�:[$�p���y쓣<��bmi ��������?�m�-O+�T�X�������u�2�xs`p?@�C �c��B�R�m`��0<ˏs,O�V�x�$�C����c�'V��[S-��K3�k?>�Q#ǧh��8~qnC6�������\K2�L�h��X��ꇶ�˓�C��Z�ִ-��@�Z�E�Y�v�5��1�ָ+��-��ָ����%��E�s��&��s/��� �mqwb�X�����|a�~ds�g{�B�DA{Q�Sqc������D�]���Z��,�)��y�X�O�-��<�շ$׏�i5��ʡ`,\�87�Z���n��`j�\�N��.��o���E�����{�ID�$6��!�?/"6{���a0Y�*�v��_:��ء���~�.��۠f��a�c���B5�:��ڶd� m��V�d������/��R�й	�����/P[uC걣���\Ǣ�H6�e�ϫ�J�PuףF�(#Fk�l��� ca��/x�����&�=��r���3�!uQ���{����J�>Q�ġz�h���I_+�1�L���C
�A�h��C��\m�&�O�j��P'�uE��)��a���������˾�ޡ��r��SbƢQ2�1S��ݐs�;n��D�m�Nw2G�Y�!ayO�O����dY,C~U��!z[��K�����p�<ۋ�|ܯ+��0�gϨ��m�az�	���5�{�RMY� �$�lz`tr0�f�� �G�v�V����:�_���Ƚ]�wC
������r��T^n�Q'���n-�xM�$�����q>!^�h9Q��c�@nא
�Ճl�n�_D�/�����g�k�a�2b��b\�4� �?�e�N맃E�D+����0�j3F��
vz�A*_���p�\�y�;o2nt��.x�9�qAa���}�1��J��
u����$��&ɾ?q�h���}Mؔ���2�����۬$j�_�[��A(�;,��+��I�7��A�Y��m���++�O��,�$�d�����ȡUFH��(�S��:U���w������!0��FͻL�5�=�g��vx^_�Jv���>e�b��Lg�V<=_�8��h��>y�0���61���j�O_��������@�X�p�:I�2�qm�/�}��RT`z7���[�a��V�bSL6��ˆҷ8��7�WUH�]t�PI��)c�1ùw}`��[��9j�:@����1h����[3d�����{"4c2/n�j��;�aw�L,a�p�`����y��C��c�kT$y��3�����8�:jR��e�	��g����`t9
׵=T��
H�w⨟(3֧��������Ĵ�1�Q&�m������߁sHw�7��1�	mK�m^����Z��rA�y��+H�b��j,NO�n�"Į�HJ����s�d��!}/��6�Š_@u��4 ��w��(μ�4��Ѻ�#*���t,0vRd�8ǗC7!�v��>�S7�ǤʑA\I�3?Y���H��U�y�&�v� ʴ�i[bp����;�E:��:Z#&��a�ua�W1ߒ��HUY����ˁb��D8�_��W��e�����eGL8_%���ȉ1�$oWu;B
�?�a��tT���Xm���ޮ��:K�pg�����$̺�w���!��vz<�:KΎE+��j����qj�}J;J8Y�r����B��t��:BS߼��?_�Jt�vMtGF,�*,C�p�G$]�	)���ȵH�͟�O����!KOz�ۤ�Wwzn_)W?(�OG��>-I{�N�)U:�a���;i�l�jw^�/�VCA�]��%�W�g ��/ӟB3��7`DsL�$9�U���er���4`փ1&��Q旗�<$�1�3��`.\e(��:��*���C���3��ѧ���"����N���=؍��%κ��
+R��8��čA�.���2�p8�Zo��tO�v�h. =X��	;�^X������`��G��v�����e�3&F@1���`�������A��;D��0m$�0������/�z�}��&���60յ�� o�v�O�*%�A��ݳ�bz��K�v^a#e2h�8j�O��`+��9�v����O�&� ���T� oA��&G 7;����ϒ�H���ə�Ab_@̏�h����J���/�R 4lg>����Xкщ���̋0KV���.�b�����OF/z��B�]��#v^��1�3�8N�N���i^������xЭ2��dE�+�v����@ƨ�(����H����L>����g9W�1�=��i�Ϯ��o�-M2��L�+uw�6bGj�� ���g!�۽���N�����#��h���!Q�!��w:'�ea��Gb�YP<���W���<���j'���@��c\��uŚ_ND(_�y�[&�O�b֯��p�9���-���´�1�7`�]'x"Rv"P�N(,�d�%��,9 ����(G �XM3�\�����H�;X���Z�ť����>l�W���y���?+͇^��)χ��?y�9}e�yZ�X��$��c�i� �S��Mi�}6~�A�)�����qh����!I)���	�1���9,L�<lL�@"��8�~Q� )vdd�*��2k�Aɀ�p��H��SG�����!���p�M�1��Q,SHCl�P��x��^�tG��_�6��5Ka�b��`� d���/���y�L
,P���0X��N�K�bg�u�B��Ǝ��D�������G�Mc+݅����8#�o�&�25D������jV~b�u�3?y��������$kY��y(��G�01����u���hA�0~l�����ql�ߤMݑ9��2$"�s�h�]N?���D���Z�#��������D��k�:�8j�yۏm��([y�d������]��z�����ioxԐ��D�6/aj�Dk�� �_f�/SFM���l��s	�ߐ�C	�C��v����V���2��5��S�|�����XX5tNGŮ��SE �O[mC5=����	1�n�G&�ô�{���WN� ����'$���o)?�QXH82y���g_k��+��vG�������߂{�=-/���fk<>�d�Obnn!_}����o��r���-�rl�����d��p[O
���kz�����P�W�/\�-�=~��4r�=��_������?�|y�TJb.��H�p�)k�z���i� �=Pأ�l�f�����(ͷ��)p�?j���{��۰<�j����ϡ��צ�g0������\��
� �|��a�b0��\�;,ƕ��8�s��'7��szr�ߞ�M6��>*�6� B��<��9i�N�}��u�	�%�ﮦ���%Cs���$�Qҧ��jm(&Ց�L٩fl=l���8��;ҾlMi����W�M���E+�zp���� �?2��摕2�����[-�Ӯ�_����B�{���W]}����E�H��e{���k��>5]�i�W*>��H�P��ݭ�G)TD>c��R*�����#�ɐ�~A�Wr�͸�x�_t���T4�/�׈v�����Ԁ)7�Lo唏8-"?Xͩ����o���k�w�'�y$2�����,�����Z�b�ٌ%ņ:��s�N�g�)Ƒ����(1�M��ɘ���Z�q�q�EA��{�a�}Y��S>�+}ͷTB�(��T��"�&�Ά��}6��>�}�;�JH}�[{�(�ϣ���%���[��!v�j��(��Y��__t?��;Xȱ"wp�+���3����kֶ0Bm�0����1���q2���@�����I��g3�"�^�NTŝ��������0ب���U�0D���7���aK�F�罹����g�+5j^��q=|;G�= -{�BY"͜B�ή%�,����^��o�l��I��HF2��-1˭�]����=�o����}D}7�����a�߹D0�WЍ�0ą��%F�9�2�$�ך�:h|%�y2������rYHJ����ڌ�)�鄲�|)c�쳻6�8'p!q[V׃=E�;L��K�Hi����Y�G���:��[^G#Z!)���Z�@8lE �^��r��ݼ�C��4}U@#H��*���Щ���W �"H���v+`�T"���/�3���8H D���p���ri�-h����A�� ��4<�X���k�0���u��A�]�<>J�����3ag'2��� �����V>����߯��m�&)�Q�H��r�L��� �g��;=�РS,S^��8Sg�u�G&B
 ��o�d[^�=�+�[z =��{���e�ο�Wj��fa%�>���ɴ��ڜ��i�*zC���Þ�x���Y�o�75&����];�:�
�ŵ.MS<�ͻ��5Lh��M�vi>N��ﲽ J��O�+[�¢θ�*�7�z���yv�%��a����Ӝ�P��Ϻؔ5����~��MDɽ!� ��0����~li���u	Z�AmȀ�sV_���q^���O����N��J3���#��m�؊2�!���FA�n>��N���df�)|z�<�>>��$��"rO���M%���&s���32�1�=Ј�����Os׿���v�ushD4�x<����H����:������-m�S-/M�/I�
�szq���f�@�M��X���bczg^C�:��/�����ʮ�]�f��0����U�	vmCѼU���D�U�� �v�2~��O�ē��ǡ��.���(銎�����hкL�_�U�်�G����^Q�O��(�pT�����]rf�	��Y�)CG���\�MON�&��U�Q=��ݯ_�C���>�.�p5)=�98X}N�󮺺z��R�vF�nC���U�lՀk��I��p�u7�u� ���FS_V�!Ô��so>==ݰ�Z��9��E����b�F��<�%���Q�W�W���f֝NlRް�E��.��ux����o�ᝨ�E-���o8-� ���t"~?���jDJ�D�qU����'������+���#0�3ٜ��zz޼'ѯ�|_�H��uN�������T���kB�(�PiӕCU��3)_ߺ��^��93���X����ٳ˞�����4�k�}����!ct�����1]�/6�a)��R��~�ʸw`��x���'/���.�����xe�n�miӓ�'999Y�$����7�/!6������N��8� !��̤�%�u�����y^�6��YNWE� v������jЎS8���dwGxCPl�Ӿ�˖����̳�u��8�3�[y��Ŵ�͛|��G�$��W�X��,�����ҥc�G�ʌѱ$F��F��,���ʙx�!36�D��gm>�t>���~��bFb)Ԇ}�kY����H +K�ԇ?���@%�@������D����-h��E�>��psE���"1ؒ��v+�����	�,�_`��/М!��h[5W�=x~��	�Oќ$��l�9�:"�Exl\���^���kV���o��l��:���y��8�G搯���3�9� U>W�٘�'#�>/>I��2��{>T��I��!�aBV�c�}��|�PݯIG�Q�Hk��Ʃx���=����h��������Q޷N�m�i�}���~��Ec5��ƍ��"R�?�˶����uO5�@li�4��oyL�Dʦ�vJK����9nF�[��{e)ڕ��������Y��3q]ۺN���͹�WD��
����X��̺W����լ�
�{�����+����3�cqM�b�q�[�o�}B��Ç�}N�&b�����7�Ż��8�+J@+��g�� l�s<�}y�=�Ϸf*�;:�<1�~?�*�)��$��,��(l��P=6�<n�kk��<	.
G}+�=�Μa}L�]���ށd1�!��n�>̪�s���>o��2h$MD���Dj�׾)	�k��o��?)�$Bd-�?ݢWg@b.�t�|�!:�t�	t*��L��s���Q��$f�79��&B��$&�4�6*�uZp*^`�M��)��aa�	�Esqǟ���β�J�vp�T!o��#�'h!����ğ�$��]���М��"?��-��k9`���q�����BeG�K+_(��8�����cxY>��1�O���Op ٘�W�b�PS���Vz����U�oj��uU�.�c4���sw{.ތN	��m$]����r�~�z�L����|�uM�e��u*��<O������L��11�H�3A�mUcz���HʎH����co��m�8�3��.�>{i��/�p���7��Կ�DL]�EtP]]$i���Pl`ĂA�u�����ԗOE\OJ\r�nN�byZB����\����Z��CS��sKh��9l���3�^jn�?�\���,#�Dz�#��Z`�'nPBI�S�K�'dRo�l��j`I-X�j�7�3>�[_ooR�n"ayI~.�%�����RNhe�3$@`�O�k�Z4/r gyt%Dr�Wf���׻(�,�VMryqE�&�}�{(����	����' B��^\��{8YH�[�$_Hf�{?��c�R�kL������0�F'��s������NIF���\{�����<�˖}�s��U��)W�<-��#��&@�$G(��܍��DP�B[��<��@J]{��T�B����ڢ�#83�镴U�tٷ��"ü�h�ZyCv=fӈ�5M���hő�ˋ���mӋ���/:uޓ+"2��PP6[ͅc[8�e�����>�~�������δ>>ӢEP2��|�7�w�k�
�}ө�y�p,���S�<����R��ܛj������w��_�T�B6�tH鷿[�XEx_\yų%UN��]� guv�_���4C��φ��o��Lm��U�)�@�D��d+x%������b��"@�lv�����IR�;d��!���^�����In�B��4i��S�6w3���x#����U�OTG0�Wწ��;88H�U.(U��k��搸�Ǟ�����l���k��sY؄@�1�*�J�R��^�"�/���2��:����5��p؇�M;(kH�������d^���/b0ݙs?Z<�Ry- ���������Ч�����Qw��Q���ޙV����I5$������+�%g�S�b���n��~�qe�(淞�*�ȗ,��!;R�ҿێȕHl206�XX 8Q���1��c�T5nӡ���ȦR�*��SӔj����:0����hI��2$K��$�N���>t��)��Sq����۷��={��u�q�)��~��%������=1��)�I��xS� G�-�?��pN��Ԗ�����4���,
��-�r�1=u�g���lC�}��E�u�ԃ�G7��i27��cҎ�{��Y���Q��&̚kW��ێ)�4]��E�{`Z=ǖ�{�7�NI��X2�·��D��t<H����%v�~�^�����S������ �X�v!4�T����c�#���4�-c�j��3�ʗ�bO֯<.��dT�DW�h�ة2��Ə
g�����=|��|�����l��|Y111A���n{�B�ȱc����Wz1b��j&��"H������,մ��`���Q���6B
�t���Kk;K#'9x}�Ћ�/�M�t��/��I�N	��xC&�Aȼ䪲��zZ��Vr��7����u�h��n����(������G���z=ο8geulnn��W]�>���422b`d���+27�,��I�5�-��8��[��K�8z�͹�-Ȱ��+�w�mS��l>ϣ*G]���-LNM��l�����L��Ż�����}�J�Q�n���:�d8j(�C�c��P����-��-=�% ���<YAJ�t7�݇V|��V{���߄)=�5 ���[8���|����]��G��Y���@���'�kJ��텅���r�t�(��[�| �
��:}j=��e��$�;��g&ք�[��?*
Cph�UK�UK�j.㯜��b֎r�7���}!Dp��
�R6O7�M�k �b�Z��9���1�{1��	���@*gخ
Π���3�}�iڔ����h/ |`S�,�o��L(][v��;8�J.�e�ށ��1_;�1��f�F��6Θ#����&�氯^�����t\#�qQ�|�8���Z�.������R.?�vY,V�7M�d|��S�5�C�M2^cb0���Gu_����d�Ӈ��F"�bccn�K|���_��f�U�V%E4�M�� �"��$������6VI1���|w�Zk��`Ւ ��Ix�F�#�}���m竾wa\����ڃ޵�y�!���dn �-�ڴ����@��=�p��al�n�������O��R(NO����[���=
m,SM�>���ܯ���.Z׍��:<q)o$�8�PTW_m?2��j'�y:;;�}�c���7_(o�z}2gI��s��Z�ZK�|�"�|(�^:�to�+�LK�?��tlJ�)0*<�l�eڻ�y�Xd�35Y�J~Rc� ��~Z�U��(o4lA5���\��G��)��$cX
!�����W���z���͑�G�U�%e����[+�ؔ%�.�}��X������VO�-�N6Q$�=�0�Qݩ��乸��;������� ���@TҨPu]к%vU�e s�I�p?�7Y&�*%��fL8 �e�^�6�����o�2��=I�Mxw<�7&��{��8Bҕ���^4�����<���/F3�8[;i��t�8k��P���P�K�����-����ص�<׿V�;{��; ��y^�՛�Gss	�U��MdM0�{����u�|��<�;v>�=�Wy��,����oyY[�n1uݼ�v�Y��	`��uCa�:R e�t��X�M���\Ȗw1�&6���[�����|fT)�JV��z�6΅��̱���%_��\���s�Yw�$����sz�������;R�UKi{� ���4Dt'����� ;(���*# ������FMf��o�z�0=���wz���}x��`���w[�|��xOrƥ������0��5s��D�1���rϦ����8��zR�⍺=���~f���[��� 5Wx���Ytmk)A���wK>���V3W�O|f$L�XD[9�������{��l^uҋT�Ƚ�CH���k�B؈Ɂ��.A��L�>bhH�Xl��]��ݟyް��D��O�(�^�Y��~�]���c���֯��%��e ����{翼Ɉ�/FQm5����'�$�``���1�ɽ��|�,�t�@������9�\g���h[� ��d���3k�yJ��D�"N���u��$+ל�T���LF��I3	�Ћ2\\�{i-ۣ��9��7�	��-ة�����t�q�ri
]�"A�ȹ&�c���`���`胭#=��O���T�=���0����M��#:)dǰ[���#�V�T>a~�Ź�#��m�)�	�{-O�ݬl�!�0��R,�N���ʙ+��`��w;t��.[���ϯ�h*(���((�}rr2tI�*�@̯�����JG};�����>�M#\�s�p��m��7 �-}?��vgؽFtm���D�쒋�3��ߢ*�Gt�����g�}��_��lՃ�=��Z�.��}�ֆ+����ߏ��mgv����7F�\H�@���n�{-05�N���I<��D�q8�7چj��r���1�9tD�s@��@�����q��SXӧ�i�H?+�~�����T��������<�J�"sM�;Q�|��YY�#d��.`������9�����`m�*g��ܑ9�UZw}�>���][0ӽ�yW�J��ִZ�u�<jӘ�o�.I�n�y*#l�<�&�V����9�L������1���.������7j N[�S��@��myfw��J�G�@���EF#�3����w�ҋ\{��5�J)|��;��'����K5�W��4��: j������F��	�I�?�jP��I�3yb��i����=`����/�>� ����=N��`��=ϓ-�4�����g먬��43�8ywA�뵳o��C��g@��� ��5ꔼK����8��qV�����o߾������>D5t�����R�e�Z����3���kI�sW��Ԛ�m\S`�Oف�(���1qq�CFY;t?ۖh�-����	B6q�ޑ��˨�vZ����S�G�� 3�TVF,�r:�1Q�������]����O��X�,�,�o��aٮ�ȇ����V�5]^�1q���!2=��S�<�z��m��jz����>��~� �G�qh>�u���}�j8�q	��2Qb��x�����^�c	�f\�&���lPI~!)O��m�~lW�KL��� d����g���\�����Mw��Qr,z�j���5�X�QAAvʿi.u�H���+)��� (J��CL��h�摊��59���S�@��000������]�wo��^�=���<�0�4hF�U�IѶ��n�6-�?��8��W�_7���D"l>��z_���XZZ�q�gb�y������=�v�c�Ho�J)%��9��$�?~�/�XDƮ�X9}�	�]@����.�����xY����r-[�eB�d�ۍ_��+F��]N:q"���o������ֲz�a��?�����Mֲ���U%�M���t�*!H<���ag�  A���ޒSS�ǚ�Xᣇ�lu!�.��N�*$5OQ�J�V8>�es����v�j��< �E8/9LA��-��>V!��M�~��߻v�ĵ�$��rv�r��$ Odyy9hy#̗�/NF�������Ϯ|��t�3 J<"�f竾�	�a��+1 {��oY?�$��$�Ν/u|�����U����}��0�����׾���u);U�%�)*::L�~�ڞ�Jw�zj?��Xc��p����S��9oo9�ȰT�|��Zeo�����%�d�qL�B�w�b��sm=�:�a��JX�;ݞXz�3{#�Zs::: *|F?�>����8��7h�ug��Yڥ�#�p�ͫz��hh�=����-rh�:����wU.~qcmMp��8�E�D]�А���m�?Y��Xp��M@C�p/�cmPd��-;-�bd�Y��rH���+��[��R8d�g��YB��$[8[�&�~�2�xN��x��N�<�ԇ�C��{}y�, t��ݞ��"�HK���嘪�h�{��?R��>>O��U���LLL@n  ZsL����I�N���J`�VI��u|����ś�}��|��~��3y����4}w<������HV��Q�){o�P�̮d�ۑU$:V�)#d��1�DI����>N�ؿ�����q�sw�u����9����K��۷o+�c����jxԝ���^��j���mO7�*��&Db}	A� ��'���l����Ȯ��Ȇ�_�i��9��	��.�7��H��h���R��ǌY��b@��zM4��Rʬ�S�&:�:���)��qb��O��Ƀ��>�d�r���3_4~��
���J�j
�
�7b=$��ĥ^�: ��,R-�S�9�+]6�s�0}o�h���r���g��X�+�5D@"&���)���ʎ$�����4��G��z�w��"d_�~M�r�xH"Le*���Y��[���-�Ժ�x��Kz��ri���������{.�Ba�7R�⩣u<u6���7���ɸ��No��6��0�0�<�X��MZ>�a�(
��Ȋ��2������N����P̼;�c��a�o��/��HXy)y|s���=�d��	�VU�K��X��-xWX3i C	m��i$	PW��dI�CF�F@����Y	�}�F%���:Н�*���&�m����|-�~�a�g�B �=�2}}`���M�^����0Raa�=Ț�pl��WͭF�8�ח��lh���h�Z��R�؉dg��S��]}}u�)r���e�s������6�!�M�f��ք�T��X���0.@z�`����1���0v�ҵ�2���T����j˶����SW���"N��P���S��A�k��z������;��謽��e�)��
v��$��-^",nG��TK�Dw��8ϝ��M?L<���A@*i��=1f%��%r�]W��@Zk�G
�:���F>�=K�!�J,t�.SN���:��U-��#��/:�F�n_�񵛮'N�ɱ���V1�P�Y�iW�۩��_Қ86A�\.'�=xU! ��N����g\��I���T��:�:�ם��_�#� P�e%�`���A�?Ra�3�P�- h�4d��Fg�KS�y��^j�#19��=�R���8�d� ���{^�m_��3�$�c�|�zu��7���C�*wBBT�aůݰ�21XY=NV�\�L��%Aqpi�gV���'�n�"vK�����嵵��ű�z޿��4�W~�jjf�d�l��m��7�E|��0� m<<*l�h#�,�kkS������E��ݱ�P�nn������7�sQ�(��Z�ݥ�\�TV����Ѕ���((*���<j�a߲l�p3|
4�ň������=&��yyy_fY�9>����<<��9kSO�|i�%�����w�G�K_;��f�L)b���Z-������c"bq��e�Qܐ]�-�!����ֹ�L�α:�%k
�O�kg��K��XX@�O�\�=8hȚ7|�R�htՌ�H�)����w=}(�G�>�V�;A�����w����bꕦ�����K[A���s��!?ޤ��)Y-H�l/w)=F��B��k�����;=�cn����N@���
�̋_jkISk%�Y�ѹ���7Qi���:1���Η��T<?{E���U����٢��v����Dh� ��oݙ�+�T<�������BXbB<@#�LG�$
�|�yt��8��j?1�e|Z@��~����CK�Zh���t_jl���т���[5u=0 �����h�usVK˭1s�5g��x���c�����\�2�ՒH�������w������^��~���X�������TknPbecc�l#v�a��$��7���1�� A%����C<^���	X����\dGG��u=��M{��^�&_�yQ��y�e�`ޥ���qmZ_Ta��zp��2��{s���A=��Y����%���Ö�/NB󌽩�i�K�&�P�Y�3ƹ���4�C1�W�!2�ٚ�T�K-;��x�qq��x���Qw�4������hσT/��@�G�8rz#K���qo���o��A��8���{�v�LF�"�'����]Avtv�J���y����.��H���x���(٢�M%�[�F��E���$+5�΅��kK-h&��V|�����+�R_m�i�)Nω���(̉����>>�<0 ��ׁ��P�(_���rTn�9�J2�IDs1��'6A�N���iLqޫׯ����B��z֝���.��7@��݋���x-y<<�D�kg�Z�}UUb��	�k�����	8�V\H��OLgI5hb�L�Qw`�j���P0�6��c$��7[���Ν?��l�����-%6�8�I�a��	,'[��h���\����/r�ξY����^�SZ_���+�+�D�ٲ�$�K������3��:D���k���?���g{.M���z0&���rO_��$�A+�������)���h�1��0ڲ�G8�n�@����!CP�P( #��R�=��b���y\S9^�~�b�Y��߁&T'�|�G�,z�I�f��Y(��v-��������u��g�4�C���Z��r"��g� �W�V�N���Ъ:��gF�-�~�8��;����z���Jի�ݻv�͠�;���k��H�1��~�{
�p����h���[�-��tQ�w���R��?���vv��|�6Q,�ÿ�����D�7�:w�}��͸흢p�K 
��G�ݎc���4W�t�=���w�Q�P����
���X����ͯ��s8X��B��>�F�����jdC�eb�\]4�ąN��/��Y��`*�s���m�EqR�R��2��f�(4�U\���	P�����x��GQ�
E�m�]D�=��ڀؽ���'i�+��tޙ���ӌ�;��TKK}�����\��gJ��\ZhGy��mv��S�jyd Sd��C�~��!%������.V)��HJ��F�����<.H��z������7��s�^�*�G 9/D���lv<�.�龹�~w���=z���6���%=B����0ۅ��Ҏ��{@��j��慆Z�Ǯ����j�v
Vy׹�>'��5x�EZ�	k�����ޘ�{�T��9���K �G�L�՟RY�
�D4z*4X��xj�5(����7Co��Ih�JN�o��*�����_� ~�R=�e<,�,݃'v`�LB��9����,���-��M���qj ^�~�/������S����?y;J������=&�me�
+������s��k�4�j�f���=������T��t����??���.Pϼ��ԏsZ�b��=��T�՛pZ����*�>��j��܂H�FMo�/��I,j�B�D���"̓BִY���yd�ʛ!ĩ�9���C������cT����⧶8#&�r�P������ڰS�-Y\s�O5q����Ai��$���jn�0�bTl�����ϩ��v��+�nn��3z��/���r-�6ȸ���}�x����꡻�����nMMM�-k���U�<@D��|�r�2w�!lܜS-f;E'����y@���:�R���q��ϯzt�B	L�i&&��8Y��^�]�T'p��^�z��$t��J�=X[�s; ���H�����F'5��B��Ȳ���S�Uq��P�\N�Q٥�TǗ�[������>y�����~��,�������2�wr��/Ma�9_�[���|P�X8-B:lF��_[�ia)'�IVZ��v�nms���� �7��/���2�y@�VTTdV�����s��bU�M��]��c!nݔ �E��5I�^z�R�K�.b��TC"��R+ɺL_]�h�z�+m�w���3���������9 ��9�o�d��+��� �쐏�����D-����G�N�k�V�P��~� K�p��`��l^0ٞ���%i��l�Q���Q�Yyi���mMf��{yAA���w�R�4i��bg�����n��)��q�����-е}'�I�aJ���昹k]��\4B��-�x��ew��?o�w"B쮉	'H�'@m�y�&m�l����~\!�V�������=Y(;w7&��D`Y�T4֎�Dc����!}[Wr���,�>O����ɣs�S���(���ۦȦ>#��:Ew�~�y��g��jڼl"27r\�󗏿*�6.��p?�"��(�,�[�6�d=���P������h4pN��!�y�����-��,�L��`�6�_�֋f��r
��Y�*q��/���(wW4�����&�B�Ȳ0k��шL�ٿfK7�*oߦ���u���B������@�L�_�޽~:�z^l����P��59� ]F,<�C0Rzi��`,&���x"r(���L�A	�	T�5 A��f�#�M�+ܬX�v��x��y)�����X��y�yX6MJ�ib��6L�<���d��ރ�0	Z���b!;���6���ϻ5F^͟�A�GEG��U�n�	r����oR6�ƪ��LD�`>(���b��w���II�m�����鯘Ab@���s]x`�rb�^ʂ�|V~u�� L��z���V����x�Y�����V|\��NP�+sm��]00��J�E�R,AP�(�]�=4@b��&t֒Pj���8^�ؐ"K6n5��_%;��+�LA,������Ä�8A�6iF���R�K����5P�1@��3�o��݌ƙ�B)�ϐ��>Qo@�d�����{CY�+G=�[�GLAAa��حE��Rc��T}
]�VQ6 ���ߚ;�s-���y5;��{�/��E���Q��h�� $�p�f3�jk�����E����k� 9`p��:��$l@4d�is�2���X&>9w����徔1A���ǯ�#�8?�a`^K�2.�i���@ �6�p5�j�bNOM�|�9�7�P��Y��g��8�ݍꍐN/ᘻ�W�_RR��<AE�N8�l�1fn�oj�o)�c#��'���?g<}���dߠ%B�n�[���W��	�Ф�6i�,/�*w����U��/��6CEF�q�3j]\�Ҍ��ܪՕSf��`�нN�� �F�ޫl666�UC2Z��o�˛�<���ߺRµ��� tg��5��<'�I��Qq�#�`P*m����M[�X �� r�V� )�O������l�KuMM����+3=!@B�Q�S.�q�|��'R"(g�Q��i*��;��;l�K8��������g?EtТ|s-:a���K�*��xU��V�0�0���gǬ"`�и����a���ճ�E������)�,S��Iڭնxg*���?4���� �f���Sw��6�~V#Q����VM��,�vq�|t8����<%`a�X��G(�鬓��2�Ɋx��v}ح4�yt�XvO6S%�ӒJJ���[v�X����S1pC�@�K�9����୏VD#
���߾�������C�7Xl:x����9����1��/��28�u�Ctnۂ��P'[`k6�{S�hw!�h����l��YE�C��HލB�˅�3�TH�g^��cC���7���~�8�n��îJ�8�i�ޝ�$�Ey�R��,�@��y����&�����
:쪒�����qR"�^y�M&YN8����4�q͏C��]n![94�d���q5>����V����^�<B��2 ~���*��zWW�J��ZN�����p�� �����KKK�;��Vl׹a���s�YYYP�@&^�o��Ѻ�]����ޫ��=����4QWW!y�Z9��A��uS �#�R 1��o�����9����CIR�{`��f�4�l�6��R'��l�^v�Q�^E8�k���X�1Ԧ��=<,hx�ʽc���A�����P�jk�1��ڃ�A�<������{�1��*,���gs�������ttt�z�ѥ΢�9�������ſQf�[�n�黻>*@����@�����=9>�.�~��W���i7xh�흝L�*�4 �/6�Һ�0���ϗ/2�%fmEF�:��z�\��ϼ��}/n꧳�������T6�����;N 1����??h�6�.�2O-�Qy�ʃC�*F>O�|����º��K-�g�R��	9Gv|(R�2�!F�#�:��2{ՓrS��aS���I(p dr������Z�󎊊����d�kn�����72y�t!�$���1w�B���w�IF�l4�j/zӹ�����)u+h	��z�X����� �`m��/�+���g�.�R%�]�H�������ۺ���ve�i��jӏ���loKὸ���"z�L�"���A������|�H��.��1�}��Y �yݙ,2݁���4̂tvK���� A"4���%y%��v�}|4ʗb&���Qh�o7�����~ỤJ
K��A"7��#D�_ju��h*�>kʤ��[� ���ci����ԤRM/���ա��Lȕ������s 9�a� ��6���f�Loۼ�*?�Dg	�c*�I���I�_3�6�Ղ�������s��m��h6=w���u ���܇V�a���X͝x>���B����@���ܢ�����B�5�2􈑜�:�y�?�43y�/�\��<����!	d��ϫ�Nc?PXĊR���)� �O������T�׳��ӌ���+���\RbƄk�"�"(˟��K��E����eQ��I�
i�?tq�C)B�;���uo����d�O�2���LSts��ؙ*Q�E��W�?��Tf;�W: ��q��Xl}=+={$˃*;Fȝ�*S"��x��.������XkH�픗�w&�J ��x���g���f)��a$�wG��>��A��^�}�|��"#��z>�LW%���$.H���S�cFӤ����]�1�on�p�9*ZJ��6�/7:��}��HO��Q�^o����R�l�[���v)��g��6d�0vO��F�[}y�;�F��C��A�s"�l����K�v�f���{v���h���K���v�C����\�}��F�bI���f%�:�{{�
�L%Ʊ>�{�C�}|R޽{�.�E�ͬ�=�Ī��Ē��e���u-��1��nX�Q��]�h�}�؛Y��|[v!����Q�ˊ���g��:�#jN.Z����ᣒi������^�����9(ం���\��4:'�0���,�~�{��@�m'GV����׹s���?d*���q)>�2
!	�e���ܳ���A��;��Ж[���!K���᥈B=���ez~�z2~.%�y���X�������	=	~g���k'�r(y��VLH����ݠg�����d�O <�Y~J�n��W(��h���v��=�ⶎ�+�p"C`+�G�vy�k

�dn>>�Ý?~�}��5M�[�|��ș���Xrh��$�-��6H�0�4��s||��]Ĝ�_6�|?�D��5G�DV�%��&}�S�D����ZtDY�*�ߤ�x��g�T��SXk�DL�6���9p���v6�������4�$��,�-�]���E,C�(��c�J��u9Taߓ�'H*o[$��P�f�`f�{�@�B�T��NT�j��:oN7Bk0�N�	=����S�ר��[�� �X.�.�:��r�f)K����G���p����ǖ�s���|�k-�ئ���P�_�ʀ	�
?�T�}��%���Gm#��^W4�j�e� u��=��5h��h.5].�条�df��������!@���RC�$�Chjv�
�o�>��P�n��s+��3D������²��Q��!y�2��sՙ�H�TYp��LΌ�g+e���;�+#�i䨕8=I~pBz�1���Y�}��tû���G��$��z���I{zv�:��&zE��h��$���-Ռ���x5��	����
���QQЉ&ҝ�x���W=0���nԝ�ݪ����,��Ʋ<��i�#��B�����[|^ԃ�����<ЈGi:P� ��q���{�$oܨ"��l��9������(^�nrO3�hyKRA��tc��W�w*�R"��@B�EY6�Ю�N��,n��H������A�/���(�r	if�r�P�X����Zw��6�p`�j�*#	a�S�3��N�ц��X/	��?d�CʒC�no�/G-/�"��"���Z�z�$q��+��~=yv+Q�&�=�9 -��s�C����wC��0��c?�Y1��Ձh�����i�c>^Պ\#�Ta3����"3��v|oCd,+�@D�����Tn^����n����Cw�CS���Uk?Gߴ������EN�@Z�ﹲ�(�z��:u:�� �NA�js�q�F�@ΐ����Y�E����8��0����y�UiJ&III}¢���իW�!䝯�}���m�#?�$�oA��	�F��z�̴���z��(����������&���N�s����M�5j^Ck�>��]�M��;���E�~}~��m�Yh?�#�7�%�;qU����g�է!h<d���N7��u��p��,�*mCł���	E�]���'j��{7胸0p�j��8�iEI��w�E�K��Y�7v	f%)��֟a�7o� �g��"�|��Y��7^�<./_h�%����L#p�_�Y�g0�lfG��l׌+�G�{�	"��u����q�-Є6�sr|�ZX�Ub[8*{,�~Be�� 
*֞�+x�N<�xL��Jx�@�����?ڭ�qZp{�D�籋�C���/\�����NY�掣�K��x���zү�X��Ú�u���%)y��[>?j,Y+|NԮ1c�.;��������j���y �9&|~���:wkѯ_�����z�0;�Uyu��4C����٥h&�9`��xAe4�m��/?�Z�C�����tm�]�J��i�mt��{�3� �o��h9׶�Z�9��H֪��l��s��#��"Q��B3w��2Y�xH����0J�K1�����׼�ѫ�F� e��1e�����W�����.RO���G���؞SRQ�k#M ���|�s|�s��p���jzSJ���0��T�����2��ow��H���?�(�1�.p>����KX�J�!�r��D��ۑ�r�?-�l�0K1�o�*t�[��|����&_����Fq�/.��k��g�U��Z�M�������H�r������A�m�=��� �x��$+�]�
�v���XQ$�
�xLSN2Of�b�|)g�����{���ljt�������d�YI�#[%`]�:��S�F��~��p��y=9��#�n��Wh~2��
$ag����hĭv&@^�"��g����b�&bd�͖q;2����0Y���%=H�v����|�G
�a��|W+���r�>�)3.s���{��_���>f����Ĺ�K����˨L5n�*X!�Sr���y���\�7����!���ͨ5�5��}��z|<ʍ��Â��E/٠��V�%����8��"�$$��{���x;8|�8�ݕ���-Z��c?�����V���K����e��\�����bh�X�b':n��{���@�C���=O�|�G[b�0�LM[�͉�u�"��缊>\��9�q��s�1��ZI������֤4\"
G��g����,�����&1-Qu��@���;�'MTy�g㗻��:�����/�k��qo� �p~�,��N�ҕ0�G�s��q����ˣa ����
�c���}���٦6��p��Ԫ춪�]k4b�"������sR+�0��c7�������}rX:��p�.ۓ�T�w����+����ml�3�CyRW��wZ{d�E���z�����RUUU7����N������j�5��ku��u����	���)|eR;�6��f�s�˅eS6���f�����
D��+`�+2�l6��-4�J˟
��fc���H�¿�i&��߳!�db���+�=Ey#����Ua`clO>O�.�)��M4+�X�*����`v�����E*�.;�����;�ئ^(���l��������5�pE����)I��pU�;n������lpne��%*�sxW�u|`�D��xh}0J��Q?~�y4"�a�m��<��e=��j31��?j��U���_�6�0C �o���~:������-�>Xai�h?� ���*�j���b:/ܻ����~]~AA���������08��Ԛ�w�ט7�1�|��ND���	���o��s��m9?h�ݔ]8��d��F�Q��4l��ND��~V�~���x+�8�>/����
�Y]	��V�֍x���Ǚ�~��,g䊗��8sN�r��F�����$:Cs��n���N�G��S�����r羱	��H�WWW�=�	����)�f�k	���Lr^Ц%U_1�F'���s[q5��P���|�O�һ[�xP�a�C��Bȵ0_#��Ȍ$^qm��S����o?�p2 ۮ^�[};�կa2m<��y�hi:�x%[��2RX+�}�`�`������e�a��/#V�be�Gk�^�	</�]����Y9�ؾ��{��;���DWc��B��E�C?��R�L	&�h��H��t='���РsE�PHP���4�`��8f����7��������[g�};��.����Lك��C�4�E�x��Q']D��^���lN7f)b@6s�Z�@��܎�/.kJi$x[�/&GR�@$����߭�#<�%ݭi�t�E�R��@��@�dĊґ�;/Q�S�����!L~�c�l�8N�z9� :"�R�-�W���I�ȷ�("��[��BBq6�A�@G���j~����~Z���-E�]��79�o��_��c
�t,
��fV�8�>�4���9��o"?�:Z5�l�������{\��?�"c��Z�I��6�ZS���R�ڃ��5�!-��O��;��T�Q�f��P��M���ڳ�拶��^P7�$H#����z�_�X�6�!c�ea"�H��A�w2QW��G )G3l݇(	�Z�X	��|��V��=��d��q��XP���gk���r�΄(�Z��?b4*�_��$�֮��U����I��-�8�#���:��N��u�=��}\4F ׬�Ѽ� ���П|���g$������/�:Uc��%���-���e�v���5Z�lJk�X'8r����^��Z;!�����N����l���42���1AQ-4�ט�\���O����d�h,����+��D��\'�#�����n���(�Rcx0l~b�1�6:׻x�0�Z&p�t�>-I����{���:^�Ȱ��JD9��5]�D�Xo���ײ��Ƽ�:b5����I��{�ܦy	��T�����������V<ؼ��$���3��rW;��ɔ��̥���R���5w�4�hDz�gGCI|�m'��[[{�b�+��22�q��?����n�O>>�Q��3��G�;5$�z�ދ:��WyZ��8�lA{�M���ɏy�w�����-]/� 'h�/�[�o^����4F$ �^Gn��`�u#�ZkS���_��Ϩ=�Qjڞ��mGVh�f�]6?�kI�N5����l�E�M�����=ڏD~%G�H��3*�ݺӤ�"�I`��'k�����GݾM[kC$�]����??�#�����ǚ%�rR}��)2���i��۫'0�r���q�ޟv���#{<������C��FC�돣�d�;��|��7P���oV�X�f�A��#Y�ץ�rD�-L�?y�PT���7F����7���R��/�x*R՜[��O�0��g9HY������*������"�9)����T����כ���BI��ͨǄ���F�'vɿ���04�m���:h#F�d��"�O)$`b�MI1��*�/L�0l]�������w=����]��*R�A����e;����Va*�@�`n�!\��%S�l o���0~�'�\ �v�n���	M6��t�U1}�қ�7OR3�S�4�v3��?a�c�y;{~�B��j{�Wn��ã��s�{H�u���PAm�_���ٽ����8�Yrd�ng��ApwJ~���fsZidܲy�)��\�E�a��dl0�4R�tE,�4ƚ�0�x�E>�>��wK*)5�-���K1w}���EҚV�k���LK~rzo��,f�[��9�Vd�ћ�☆\��G;�?$Pj���hT����R�c�z�D��a�u|����M u��=�]����?�0 $U�h��N���~�%�[KU'���L^Q��% ����+�ϯ+`��pho֚��_��fG#L�luv�sc-P�+H�Σ���g��ϫ��	
�#��4aUKWD"O��ޛ<m��3�U��	��Af���2P���Ғ��E�~��Z ����hī�xω����=/3��6X�WO_ެ�� ��Q�8�e/�F�D8�=��c�J��N��TOꆞ''(�D}��R��"��r� ��w儜�F��Z���mRC��/��t�2��T@�`��˻e�9��@N^��K�.z:�V�Fj>�6w>5x8�S�k�Ba�t��G�2FD#��Za�>�L����s-qF�sa�?H�%K�wM�6�Y������	���.-t��>=�iR�C,f��wc���wt�UO��9M�t)LR̓m3����+l/S	�<6�s��)>������{�\���Aq�_�7EAS;ܱ���WL$ztC�?���ID�+��!�+�bHV��N!�LdIp��Ǭ1j T���#ԯ���6����_.g4[��4}#i�v�ߞ=�&%+t�Aώ�I	�2N����'�[����R+���;���h�X��;�[^5���Z	�M�mMM��P�Z������� ��9 ����������Q%���|}�ǀ�c?i����lNg:�ɳ*�~��0bc��lVE�l��l �B�[�'H+_5�'�.��B�����[7�kEH����K�}�t����؝��Ȥ Qc`~�7�E?��IYy�� �ֻ�5ZaCK�t��i�`�gv�N}kkk]Ss�N���{�Zu��N�*+^5f�Msh�g�|8����M�2��_=e!�;���ɸlv�7��_��v��M�(|�6k�X�2����n/*� #���eT:k�"�wp�p�'VM�6����0�J���۵�]%2/�&�^�:E6��E��T�#�]F�{�1fi�@:����>�vU9������jqϲZ�/���<������h�qq����n��%rM�j�۪ ������88-S���C�D��j���T@��sJ�7�O���,0҇��!����zP���rр�٤{��l�ھ�T;�T�!:��/�<J��&��i��-T�r*?~�W;RoN�Z۞^`�4fd�[�N#����1H��/�g�qթ�9Ȥ� �L�&ZP�\������#����5�:�o.�&��4�$�ioQT�X��B�¤��~=\2cgO.�*^�X��I!����S������+��ܹ�y� �ޟ/4b�n(�$š�?рiL#�ؤ���RG� pQ�8���ı/"��KG76���"l �	z�g��Эq�UV��?dX3�%��
>�>�,_c�)�}�
t����D�4)2��7zN��X���?�N&��s.!�����'���
bx'oH��6,��N��G8�(�&)��q�)~4r���qO:j�PB�i�&�L_���?���. ��d5+���t�Z���o�Qٵ�����/;��ݴoo�GG7,I��L@K�S)�֫���r�>�����������V7�\�[1R�c�z�A<mS�k��~��א8��,�,P-�7p�T|Ƕ5W]k)������PΣ�ū���\)��`��Q��=(�cNZR���p����p��! ���~L2��/��M�������Z����QjUgV�@��ٟ��"q�U�U�^�ۮ�m����B�f���|��=�-����	�M}	�.x1�{O9��L����y>ZB�R��Ô��F'�B{�
Z�v�NP�s�t������_���.ȩ�� P��#>���_�]����>��ʿ�q����/Oy@��x�4��="��_	BK5p��v#��,���h��4������=�F��S�Aۿ�p�*,�������'��p��#�H%AowS>�r5B��L������z�W����gg�e 
��s{���r��Kk�����HV՞K:>�Iz\�������wYY�c.��G�������]��)&���T�9N8!��/R?�H��17tK�+�1�5�.�Oc�E�Yr-�',��Ts�����C`���nl��C�~]Sk&p��c?�Z:Dp���U!��ۇ�8H9��x�c����%i7F��d�<�ڹ�Y|�0迎D7hu���,},�@�_����%�!l(A,zz�(Tm�b ��5@��Y2�bx��4�"fMi����)�,B������`�|��ޞ���(��� z�8m�F�{̭��vOi;z�����Z�.:�z!��R#����o�������JO�s-�n0�Թ�C��}�y��9!�g8�+������dwVmuꯜ�q��jsq�qs����X2�{8@�5z��Ub8.J�!1W�B��"z=-R"+}�]Г�V���q��A QVv��ڪM�@
VH6��,*�KO�8䴳(�^
��XU�r`}4��ϫK�__��Ъ�ӿJ�:���^�p���:�
�?g.
�}��þ�~�)�_�	�V�QٰcG V�*� ���T�2�F$,�>H�h�Ӏ`v W�]��l�]�
��m@r��m��hzJm��#\�����S<g��/z��[��H������ɺ�LE_J����|�g��ƌ�A7�ھ��V�g�Nו��� �ˬ�t�WЦm�3l&�)]�h���t�3�D+}���%�gM�f�]q���j?�~�ދȣ�cX��8��w�n�PfPt�|��%�sy�:�N	����"ܻ�L�S�#pԜ��އ5�,�O�O� FH����T�[��
����	P��I����$��T���x@嚕����ӧ���z�'�Z�&��~�z0a��t@�9[�%G��Q���r���b!��D�-[Q`���'4~ld�S}_��L`��<�����[��a�W�Ŧ��Οģ/ځNh��Z�p(X|1��8s�Zx �-�A�x�ʝ1o�t�ʿ[��\C�ҩ�\� r�K�hPuu�������eĩFDB��R	N����,� �\�}O@���������"�F����O��.E3��pG��)��s��Ȅ��P��Or�\�3ۀ�g	d�[�Ag���U�hE�����R|I>�~ŵ	�߸��ٲ��7n�5���fd��X���O���D{���5\�G �klBp��Mv ���r��? ��C��(�J����)d����BP)�U�y�C 7F(�����g(ݨBN��=�ѹK{�5�7S�g6�_7��~�rp�J�f� ATj��
%7,IK����Veh�r�a��<�p����d{�d{���/�M��c��m�~ ; tE�tp�돣N[�p�u���a,ep��	��t~Z|������I1�s��������\d,�N�HZ��W6묆d&r�HhѤX�|T�/��vPk'lS�?���	l�K�"�X$P�c�%RtM�&��c�W�8�ٔA��$Z�Y%����4��	[^�]L����Ԇ��џ�vw_sQ�����y'{���^�.fp�Ŕ�"6�}�liX���j���v�+����8H]͂Y��>����ĢTiJ��	���g)6)}�B+�߿ �04-^ı,BO#I�PPP��ugUh����r�t�y�/-���h���l�ٸ������3�3ᵅ�a�d۷��h�;:�2Z}��aq<sXq��귌�?��Je�`���M�vI�B%�M./;L�mM��7`3������5~������f�͚0�g="��4ʧ\Dr[��Y�[��O�ݹ�˴�P;����_��>��RO�ٔ�bX�� �*�=��p��p|��'�k�'P���̾{ �6����ݻw�0��U�[;��{�㘋~وA܆����m���ǽl.cT�c�@��.ES��9wk��g�2K�d���J��Q�z��!,jR�_GA��;��;UJ
 
��ƈR.]��?�g��/S���A��C�#Nd�Olx v���a�h$�����_�H«(*���Ř�K���D�-L��{�b�[>D�ӝN��a=��F"���^&$���C,0�կ�����[���/��V5��T_o�����FĿ�8�� &�@��bPw[�������i��eh�A�4�N���T������}[�tS��Ѩ��x�Ъ�e!�<rؒ����E��'3����ǧ<�%�/>�p��]iz��7M�1~v{r΢���И��Ŕ\�����lU�����B#9fn���s+������tz?(���p��`�3�n^�]�Oүç��=L��?�خ!(`�=\j�I����A��)�ޚA !�X�eZȾt��1aͰb�S�ܠ�3�zI(�ԓ�仢���:5h���J�$�(H9G����HX�g�434�A�,lk�*�5|?�"��<ʬQP�y{���$��45���3Yvf X2����Z]B>��~l}��p�	J��-Κ�'P@
B$�rn�y���Y��~[;�����~���y�̃׬��rJ"gb��D�9+����KY�_(��V��ڔ�.R].�.�Z!8���ݘ��`C�S�z)���>��ٽ�%?��jn8AD���״���-]�ZX���~. *m�NS*��,za�O.��&h���W ̣������R˚�L�u��oA�Nc�� �K�M�/�O����64yL���n�.[�D2ڬ�͈���S�j� ��y<w���)��}�.������=҄$D�Rd�ԉ"߼L6����c���|!��\�費A�4�rڎ-�Ct,�ct�y �k���R!cT�|��蟶��E���XR$��@R
�#έw�.���E\#���4gbv*.z�Rc�T7홏��I�د#nt�����?h�=�,b3NN�l����c	6�׼M>������Q�	.���SK��x	�a<B�E.�Z�]s�Z���߈��� 1��֐�D�=S������T����V2Zf����H[���ZE��\�"ԕ�F\{��}�E�-���е�_o�����N������|�����B�T�����Z��KS���<�?�3���%K�V�A���+z�Ϥ�q.Q��':��?�ُ�=�׿��84>ZA�.&�
��Lw�!\=�3�=��'Xc�$AЙ�%����1�ָ����^���7.w�d���C�),��I.qʐ����{߯�c ��p��ҝ dj|�a�� ��B����Ʒ#��~��}gy�oqg7�C�ڌa�m͡�ÁB^y����dv�;��i4�5��]�\~!��Q����<p]žEc��>���P���c৞���4�8��̸�-����L2����f�;t+󉦔��F��l�dK����,�ݡ�c�pg�E�iR���#T�/��ۑ���fQ�)�߈g�����^6�3����!�bE~�&��ş��X�ؼOkג?�����73>�����
Z���u��{�旆!�������oP�ܦ�j��0���|)l��S'`S�P��?�S_s�p��J���9����d[�T��,�Y�Е�{�QW����<�G\��,4�i8l�A��͢��Tm4�C��3�P�$���g�CE28}��З}�tZ,�L_%�~�Qټ��]�F�cv"T_�:
5�օ٬0j��S��m( ���1���61���2�)�৮@>|�	X�[51��;XSwy�QG��\a�u�?ſà���Gg��& �f�Z�% �Sg	�`B������9Ȇ�Ш�X���7��x�d�	�n���!��o&�P.��.�ڮ���e��
��K���G�	�~V��}2*c�UC|Z��Y�����B��$��F�5 ����7x�jEct��݀�l�U$]��{���"]5�~���B]#4��acN:V��OZ֊L���ts�Fi����5���	z8�N���4��2RLD����1�u��~�����{��f���,;w������Y.��aX���bE��������F+��n]�/5�����>y�[G�z�J��f�!6/|5iv���h��Ȇhሃ�;4�#�}�������������Fb��%;��DI9��,��ڧ��v��]�,�z�)s�97 2����DLQ�dKl�U��9!HoI��ܓ��J�.����E��ܜ�[���T��{�E9�c�����W��k&�/�CշEA���=�%W����_.I�s%��~�7 \�:x\�|d�U���W����c�ey����'K�._����B���/b�����E�^O�F���"ԗ�"�� ������>��h��
]. ��ؕX�H�9�E~)z�ցb��0��&�LŹ����_2����\y*������W��������JQ��dpvr��S$�,I!���r��띾�h�&`D���&�;�i�J3����F2jcû;��Žėc	�>g�c�ZZ9��O�Ζ���5Ł(���T�|����`B�`*9�D��7
h�������1�/I�e��4(�$b2�6�k�]���:�y��@wN���B�f�ϒ�>�(a���>W�=��x����R�A�{8�3�����/�C~�4:
�8�^ӈ���}��:c3����>�"�-��ZhKЉ8+r=fj3b C3}�_����b��c�ae�Q'w�2�BefJGcP�c�m��Pz�q.t��`�%׼c_;��?�]���q���{"�wHE3�VO~(�|3�~�j����.���g�x�*��*,G7���3��q	/�Z�:� �uh9fA�Yb����@*S>F���>:<�i�X�I�-���W�����/��>׸Ys�S��7�7Ug@����h�SrJ���袅����!���>�&��M(�7>����l�^�H3z��sj��g������;��,4_p�DW'g��;Vfl�t��|_[.%�m?/d�?���8J7Tor=8@:�2(~�(�R�W� u(	���W	�Ǯ����`n\<p��B�
�-��~[㪙��s�`���]o��$7��O�v�G�<;h0��^���S�_)1���>�u����&�+��e,�R4�:�Eȓ��W
��O��$���̠,D$x|3~�~+�/ ���ac��$R.�:�
p�7�ǲn*�:�����i4Zjb��k��rJ�:�>o��R�U��hdl"�P� h= 5�k_�f��A�6TJ��	��R:4�s��ZvO���M����K��5��O��3`�X�y�y��	��I9"^�E�Կ��x�g��@,(L:��,*�n��s�$���O��$ʓ/��
���2O���=S=�BmBr�a�!Q�?�n	�٨h���������<(�x�~G��0)a���bXu1��p���"g���R '��������E#����=���**aE��O�����~6ό���׀�u&�=�и�<`�գ1����_;�)Bc�}���Э�~W�)I�O�a�,5*�*,1�1��a���_��'�I!N�Ms�f���ޙO�;v�-�p�?SL � t���U��H����\�e'O��%�H�E7��#E��H#�+�>��ܿ�cH�j4��cȴ1(�
�°�t�)z��;P@5=�H�?0y�$b>�)&�S 29��`t��`K�T�bqhss�}���F����|{N��p��r��L����L��f�:;��sB���u�����,�E����+���z,5Z�m�Q7��\��}�e�B&�0'���p��-N&�(�l����?&��āl<Q���5��c����i��w*��iSrf�wMxI��UN���W>�s��� .�"
O�d8w��er+����rJ�R)�����1¶I>�D�8�<X���:�_5IIո@����1sS|I;6�RDq�: )�,�3m�p9'x14�#���ƑOY'��!�9t�5z��5"F�!�����;����c�9M�wt�����8F��;Y6~����J9� �BY7t�+����lY�m^8�p�,��E��X�d����x�u[4�7�8�
h���"���� �{��w,,�;���r#�S61$*c��IP�

��И��q%��Q�$���`__��X��a
�M�ad&$��ᑃUd4�c��9��A���{I�;�����ѐ��$+��@������v�.����&?đ0�@�e= kj_m�����xX"t��$���bݑ^�"��������@�+%�Z�/�?mѨ�֝�&;u⡦�͔�{�=9CE ��
�Ñ�K�@�@ɻn��X��R�t4��L�zG`�ba��D�S��w!���^vݤcoBW�(3tX������Rʬ���Î�^���JGޞ<Q��s��e�9��$1I���PRTU�{d�����7�[�˷�y?Փ�|�I�XF�޹j\m!H1x_8R����&��N4��U�"`�>%�Et4X&��G����{�w[���}z�
k{]�[�{�0^/��u�[-L~B�:1�;m�\�IkO��^��@s�"�p=�*@u��'��M�˙F���C��d\�]L7	qp�}|�{��1/��'�G�CtF�ߪ�L-w�}���l��%���^J^�ey��z,N\\��|N�i�WT��Β;����B�T�e���k
���!"�P	r��vbV�yu�_�]h�%��K�m�f�����Lx\xZZR}m63`|�J-9�r�N����l�{^�9:��U����i©�'�<�c��"i�<�,`�oѦ��ﲗ�y���Nw�Hɾ�9:��}ΊH��p�H6&��54ۦ�_9"����+����t�l�x�ĭ9pp�J{�}�p^�{���J_2������/P÷�
������ ���5�!s�:!��l��'�L6s8�*=bʬh(��ur)��$O/�H[z���C�>X+�Q��gX?�E�z�^櫳���`:�38�(�r ���T4����?�P4���3a�!�K�e_��m��2ƅ\Q`{����wq#�o�������T���w���WS��(�h�QqoT�@K(1J ��&Fp���`8I[�I;i�8
L�K��~ʀj��ݻ�\WJ|�V�/����}����K� �"oh�SH����_%�Ţ�B�v����w��7��c��6�ׯ�c�F��۝"01�b���"���B���Ξ������.txoj\3��ãz�O�hB���qYG���{��(��d__�$�����ih�F�l60���U�8׸�F�!/N�PM�����G����@�o�2�<	=ᾙt�6|�8G��z8�v5&���(�ިq�⥠���N߹�&�&J����:;!����Q[7�)���(��y��

&������A��]�3@W�Og0����
���J�-$v�B3~b�2b�|��i�N����,j��ǩ�����w��0����&��L^$;��
ੑr��D���dQ�S�+ާzUu��S^�?��]�@?�Ky��*���4H�L�8�	f8[jp�B�/~������.>���b����|"���q�.�5{������^�'��	���m`��jz=���-�x�*z���۟gd?q,��#�X��(|$�p0U?��-�g���E{����er1h�?%*�H�?B�-�GS����]Q�/_�GU܆nA*����;W���Ls���!$���C9ڱ_������"O�U�H�& �?�=�_
���\�zd�A�)��㗝	��7Oz�:��׍��3�vjJ�w�z���ئ?F��kl504�e��{�W�sK%AӉ�F�ŝ��w���ûζ.�����D6[�!C)�^�1"S���L�#�`���hm�荛�Z
1bv38��B��>n�}�(q�TQaoc�+t'<��ߣy������/����:텒�Tg)h޽�p�� w�=�K��7ۗk8e�@J�"�$,�&���=�u�{�tc�7fzG?���ֱ��j٠�w���j{�Y�kO����%8*w����<GR�n��hc�n���T�/�W�^U�A�h·3�*T �TK����W?��J5���D��� _�E�{�'8v����	��&���dI9:'��As���^���(�Sm��]q	H�#�]����!�
��_���ip�B���ÝUA�v��,��~$��aa������9����_8����/ۧ�������_?�o:�|���ၽ��2?8�C����	�}x�i:[��y���0;�$��'���GSߥ�Ε�����/�w����<C)�g�*Vy�����c�gy��ˢ��dgUSc9� dB�2�۫��R�ˀ?��(E����m�V�st�uZڝ�P4������_X�N��(z�MY�sM� ]�,����$���$�����:{;�UC؞�s��e�Q)$��.�8K�7
��=47Ϡ�憊t��|��E�=?�����KZ*�=	�ޠ�s�:��l1���R����bj��T�>��C����ZJ!����]o���(��"�_�|B�ك�����G!�+f@T9�l����A��� C"��N@���9x� ����l,�����J�0��������$������w������H�{l�,�e%�L꽯8LR__ߨʈ�̚\a`9�Z���c<DBkk~����=Ѓ��s�%�=��=��M�U$�W��/�^���-��2�v��u�)�)��?�Ru^"�Ǭ'��#[�:;M]�Z��kh��������7������Z9��ٗ�De����N�'x�*��^�~a�����f~|V�+��řw]������Sg�ST�vZͬA�&әq�*�%��T�vxx�a�֏~���D���v�S�`�ꂆ=��6���_?�����W����H�h�Ba�����!���4{"ۊ�i�4~J��+en2��Ěf͋>�S3�� �j����iF�	�hP�H��-j�oZ2���1\#���N�M��l�]X���$̘���u��7����&o��]��n�^f\(~q��֘?�����ؚ��������)�UiQJ2Qq{O�0'C_�X�NO8j��1����A!
O0��A[Z�\Z͔`V�>Kj�/��(�E��bȖ����MD�S���K�Ey���b���VE~v1q���歳`�*w�oZ��Y��߼m�Pv�P"_�x�n/j�=N+�5����ϟ༸q�Gc��pt�z^�lR�,:99i����tdk'l?AA���Q{��wТ� �F�.��>t��^Ԅ0#��h�I�`���r��7F2���G����[MM\����#Y�d���|p�4t:�5P[8%�'�P&U�vC[�B�N�)&o|��&&&B�@��GB�<��Y��;�iM'$��,bo���MXCa�t�!X���0
WuA��s|L�G��Ci���^8v���Q����4���5�i�`/2���	<��SE;t�C��D�@����4�U=l��z��Аe!)Ŕ�"C���P��@��s~]M8Z��qw���o$���0a��go�׏#�s~��N$��"N�b�uH�x��CӦ�/�F�j�У-EEE���<�U��ΉY�R��;��c�����
߉���_OXoŻ��(~j��5#x���;CΜ��;¢P�9ă�2����_P��X]]���}�뇡V�o���D܍ T��|�����ih��0-��
�6ι@7��5�!Q�#5�~x���w�l��y�꟏����ە����(__��������j�%q�y,4��nTO(Yh��o���/�㷭���f��{�>ڛ*}��l^↝�h1�|���O�K_��]#))R�Ss�����}7O��,�j�/[/6p�P1;w�s�1⛶Q;��lS6޵0�?�}o`p�>�F�����N��88^>�-�[Oh��+)�k,��MD�ׇ�I�S
`�,�T��nJ��+��|yMM��DJ��j����� J������ǀ��� �O7Wr��!�8�69C�?ws��~�����&�Uό����3�/�Mĕ �i2�m�p�z��2�3�A�J�F
+�B��D)�ǿgS�e!���$�L���Ϧ�{���R�d�7p�Q��LM1M�]�:���k��#����[�܉��V��K/(�ry��`V�F�l����ki�Έ� և�D�zf��!��GM���}�!��'/��K�<�˚�A=�q�i��ё�H�:���h�14�7?m�,2/�_Z"W8���X4Λ��Ѥ�ݺ,�;�u���$��=U�L���N����7�I���V���o��af�,*H��m��q�\��ntM)c��#˕�L���w�gk�J9"�p���g�m���$Hީ�y6�  e��W^_��ӆ���*R/o�7���LS�J队���T��_�A���*�|�>e��yۗ�cT�X�
�f�o]�N��N>V֮��˗G��Iզр������(u�2*i�w�|
�R��s���P2
�f���̑Y�8��KY֛�
;}ӫ���_u%r�H#v7�-|��1���V�1��T���3�&S����-��~����[4o�zz�n�rwwO�����ո0�Omqx����~�Z;��:�Ȃϻ�ƅ�;�����I���[���5�1�R{<�9���~¬�0,<q�{� ���jd��W"F��t�2�z���^���7�*AF�k��zt赙	5I�� 
�M��'-,|h���,B�\iԱ��nuR#�͂Ỵ�-�#��8
Mu�'?�:kk?Yr���P>;�I��U��� ���a��Io>G�ڙW�5��՜�6� �N�k�h,��W�m������	xإ�2���7%��D�+a�"Qd/�;�x�3��O�c�7�O�GAՐWP��"���ق_�/�^�)�g^��!�OL4ϯ�Ȟ8��%ti�"�t�c�f��&mn�Es{�b� bK<S=� IG��jהOm֗�KZS�20���<{�:�h��(R�~��1�N.f<u=��b���)�W���_mFpݩk{��B���ua�~Gm?��n��K�t��A�I�������림j��&8�"8R�;�[�n_�L*ICS�%��~?<|������0���6���R:���qN�Hd��`�� �}�y�Gt7������D,5Y�8(�2�_[�B�W3�8���}8��|��#h�Y g����`d:KA���p��N˦��0�ε�~�6��jm1ֲ)�[k.�%Ś!�fJ��3c���tC�FFF��m� ���B�N��Rf?rd��TG����)�����M�D�H�.�s����A�qXx�Z"��ن��Q�w�ɐ~4�`�G�n�ӑ��1�~�<��Z9�|��37B���b@(;�Y��x��;������mL&��k]U��\�媦�F��s�20�����g-N�x����6�;�p��`���D���D�n������L�h6[7�Ά3�l��q>8�g�c*��J��ۚw�$>)���?������}�"�h�O��0�ą�
��N�cy�L�ΕH�� ���?@+K�|c�|�2<A���Z�G�тn�ZKu|�ds��E$�U�a��8]C+�2���p�����5���������E�sqX���7��!5��g%�{>|�.���#<��A��*-vzEO%~n|��w��i%��&���T�:�'_�A#5
Ŷ�{�����m�[.���������{�y A;�׃4�V��`�0�C�m-u��z1&rf*v�|k4?�zGcp��]����@�4��zg�\�������6�{DN�v,I�^Ki�aV�G�Ld������S^�� 5Qvt�o���+4%}=f�K�g�������7�൪p{v�%�瞱Ǭq�8�&���\o�UR����~���QƗe�[f�����RQJۺ	��S�a�JŏVIۯo4�$�)[vg����6?�Z�s�y�޿}L�!k:����o,]Vg�����<���q��ӬϰDlm~�m�J�Xm)��Q"���+w��9x�Q2��xskk/�壍huv�t0X��R�[
�>����-�a7�Q��ϴ#�h�� �k|�M�WSS�WǽX���'%���_&�.^��+���kk���>���g�d�~�鹸�FKٔ{�8�[�L��l{���47����5�yB���V�ꟗ���D�;�$t���/n7�+����9xvѩl��(�����2+��%L�џ�J�K�A�*�ڤ�_��6���=����[O�b�&��ws�m���"��M�� ��#��n	�d�:2~fN]�фh	��P���p!����j\B)���!��B���9]������O�ɚ-o����_go�Ā�	H�J�P�>I�/�q4�Q���!����Ё���ul�FU)jس��q~#�[��]�'���<mV|a��/����eW4z5���(�n٧V��T��ߴ��^�i�/�^�EG]��G���޹N�~�b�K���M�5��n�o ��7�_Mp�E$�6�c!ͅ][�n���JW��^�P�B.@9���e\� �A�6��Z�K�x���b�MsGqx�:���k����ƒ��h��
n_��`���qr�PwL�m��R�Cy
�tJS�"�ym7?r{d�t�ٻ.-@�:�����������,�7B���$��9�u����X�X�Jyn,�ߚ�1|������5#N������5KLϥ�e'�mb�t��^��Sm�۰�[���[���]�����U/�BSc<*߄��T����om�s��\dd��D�����R��=m��#�q�Z�����n+�����e�L�_�Q����dk�b��+�-����H��X�ۙ2�����ȭ�yU%����t��Qz��*��],� ?ou���^���Bn]��1h9��T��D����I׆��wC�Dlv������s��sن/J��0�fz�I�=��Ԫ��G���(TH1��)Zh#kt�R�`�4� qxtѩ���#��2��=�E<���s� `tE�>	���fӞ�y��'�΄\z�&��Z~t�+�ўX�|Q�/��l��D_Vh��X�S�i<;��l���l]��97?P���r:�C�_j@�Ve��ȅ��o��ثu���R�ᯚ6~�6=�җޫT�U��af8�����~_!.n� ѤN�S���w�8�y�m=� �rۮ�YS��:W� ��-��F�$��D�]��7N"n������`��M,�Y6Wۻ�Ԣ���sEI3����oztˆ��ԕ@����g��6��h�>�n\BiZ@}|���
����vvBs��w�#�`B�v� 4-���7%Ƣ`�����{,��V�{��rW��}2<@$o����:Ԁ�����"X���z���\�CYF�+TI:�Դ��O�����G�M�2��u8�v�|j�H��!���?�d��}�O0Fl����=:�G�}�C�){���ѐa�,MJ�Q����2�v��P=����R�����ϗ"}�L������!4��`oME�S�a�[��y*��G긮}.Fh���^桇��&���W�աz:;���K|9���#��1�k����Ҥl�>K���=����j'n���|q�/�bX�ܛ�l�QQ�۷/������tR����1�+��ܪ"��r󡎀��|�����*��٧��	�I�k=�V:��!���]p�kN a��$<�-:��r��#R(e-�gI�
�AIiiO��qO��"�:���x�!߸�ܱmm�'�˔F0�yw+(����~fy������[kZ���n�5�_:��]<<�i���哪L��.�v���\�����[*&Ĕ[���{g�An��Tp?A��W4�g�Ζ0r̋\J\B�����|���7���7����_n���O^�Z��\�L�.J
3��N���aI�;!0in�Va���{��&�����K(�0gd4��|�h:��k�K@�O�d�m��J���h����ʎ�3�l��ZӃ��WV��P5��xئ@ڙ��*v\��gN�g��1 x&�F��'��aE�Vyj�{���>5%�3�vٻ����{`�-N�)d���}꣬m]��P�i�V��<p;�񿴟|������b��usrz�3'�զZ�xH���&�ێ����V����H�����V6�w��x���S��S{j�?�ȼ�_�}Ɣ{��a��yf�M:d)v-:ￛx�Q���*Pp#J��������Q!��V���w��9O�4ϖ���1�>D�S/�����]�������H�%�>]���b��J�[Y�ۥ�sN1�����ݨ�/&0L�sy����/�^�	����*����֪}t�5�]㯉��ޱ��Ah\���ݶf+�3'�bemYEr�� ci�^tdѕ7l0D;o��vi��w��&�T��t!�p5k�K$�د���4ߕ�Ȇ��x�/*���/�����!sDg���~|���ƍ�/f�	a��^j��SiD�J��p+�^�		W��(��Pk��Ly���+[`#{6I���%U�r���R�/o�%vQ��Z/lv1��Q�`�Qv�J�hsrNj�Ϟ2�ц����y�W�c�և2,�K�;F+nʔ{�2J

��3�Hc	�R��$G�BF�n��ϓ	�AO?��.��N\ӶT�y"z?a�м���ߊo�@������~m��a&�b�����[+t�:����@���8�3�����@�#����{8��n�TJ��XbxR���?!�+nIl��1�����wG5�@��uTT��4P_��Q��r~�	�qq[����F4��Q\��ص���ke�������Ҳ!��d�6�:���1kݶu�X1�1����m�v�X��(Q��\U�p���������+Q3���y[�[V�>^HLז�.͛���֚�r�<E�F���i�=v�B|�5��k"���w�����L���Y�ؒ�z��3�{ ^��.��k(S�9O����6�S�([��,�`�]��wN�%����H>�?����|�r����6�L�R4��_h�Ҁ�DG����ǖ���C/�B��j���!���󹓓�r��/&���g�V��e@Ơ\۝�߭�{��Q���=�� �
fo�6��VL�)����K
�WU�-�d���Z��z짶���A'�-���im�#N�h��ݛl�49�`[�����0��=i2
���8z�pk����"�U%�#�d��������5��b�3�@9�V���Bm���N�e���Ύ�'ۣ�1-��=�����l��	�5�;�$5��=���c\�BSH;2�v�1&D-sz�:!Y�]�m�+)ϡ��O���ʚ�w�R����'S�U���~�sh#oߠ6�;7`����ߗ2ͤ<^8����t��H�lL��M�=�����+g���({{�ܱ�k}��3��!ʹ�΁k5�~a4}��!��₭�	d�^�_��:ў�n�$���!j�Y��#��8W��/y=��HKK;��%R�KC�]s��R��C�\�.��9�ݢ���te|/��J���=���8[ xff���X1
7_X�EL:kQ�]#$xS`�l[j�M������*べ��u�������ܱ����;&���lgV���**'C�S�_�O{~�@}eP�3QU]}6�]��v�����ѽ�I��]Z�<�'ݨ<@�`tD��KJ],�̩EO��mʕ_H�D��1U��?NG�hM]�ϱ��\�iK�Z�k��ы�ł�'�W7Co���:�`O�Ng0vvu���Zym��^�;;9U:�d�.V}�H��������d�%Q�����/�ɚX/��Y��8�W{�@�s]�K��5�8��!z���r!]	^w򍍤�Wv����O�a�������<�$�8\�=66�r�Ն�iwW`�fi��v�^�/�����iY�Js�X[g�8�������S����j�Vs�������������h(�^�Q@g/oР���e��� }=��X���й�a=���p-K�����l�z�F)��T�4?ĲdX��O��<k�r�J��>�7����o�=���0���P������J��ö�]j��?C�lM�̩�6��u�PҚR딗��d�n�91���
��eϮ���t-��?R3�S��4����G�YTm8c�N�[�)J�ν������#U�uuuМ|�guqE����b$�-	4����9�jJ2V��Crn���f4+6��>��GP`jjj��õU��?�_�h�>��㙪��k�F���p9�:�����_�ɘ���P�Q�Z��yP���N�S�hjc�ۋM^��t����맇��ˋ�/�,��c��y�,���s6��lv�9����tS�����
`e�]��(]�P����QQlH��� �U/}6ܘ�h��R�9mĘ�d��f�$���4�[i_�]_��)�tw��)��������/x%�߅��T*_O�b�V���}J�س�j@9��1�����#�2��μ��sԎ�l��4��TR �~j5hju�d���|��O4�\`�4���W����0P333#��J���eftv꽯7a�C�&4������@�QhR�6Bj2�~R�i%.&����m�p��N[��[���.���u���� p��sSRO��	`Z]�������tG�?i�����>H&zTKxn���p6(!o�_u��d���:��3���5~ȕ���P��d�i �2d�k8�~Q\]/;���iy��D��_]]��g����� ��ۗ������f���<q8��?�j^'{wgN}}#T���	4s�sV_�\�{Rô$�4Q��{���~�q=�mJ(QU��-���7>�p�a�jUԅ�Zf9=j\؟^ϻ�sK�Q�"f�\k�[���_����ƍV�L������J]G.q(ΰc�^��b�@��D�|�׹\�ܭlI剉�@!��a���gΜ��033�sT�*�� ~/�2�ATWww��pCn.�����yc�����������Y:��glH ��+*)�?{v���,�R,���L&���H�3�b�^l����zzzofX-X�̡�4��dB��v<3���(�>=5777��i��-X��ǂ�%��� �0�2c0|�~Sߓ�t����O�r����ϓ/�Fd��K�`�c��s���z@B?��z����($�A��x#G��nF�:d.� �b��J����V<��Hv&����lgCj�i`���Q˻�űB�m�#Ma��r�TjKu�\�ˍ^��s�$+�Z�A�	��ŕ�/,��1�*��xM9M��G�d��d�A�W,�5�M*��þt������8�\�З'�ي�;׶�|�������(��� tv��ܼ�����&-��?��?5��LWW��/eۮ��/�er�G�:��:- %��y/�<Ew?��j�R����ِWZZ����K��}����ǳGmI�VZ[[�Ԋ~����^=�?��Q'���={����q��{��@����su�N�]����h�$������{N�-��'R����[��ͱ'��q��<Q����Q�B���A��%����n%u��z����͹�v���\~�&ό��o���j���gS`)-��"��	�����9b>�
�OX/�Rh�UBq���3}��J'�����0���'�*  ����^��b/rC���;��/n�L��S�cf`=��Ҍ�-�M�nħ֦�~�c���O��Q }�����H����e(��q	�x��E"��R�|�
᭫���:���߫s�\���y9������(�]��*�S�+=�9�N��瀱��������a�I��{�6~�Ħ�-��Qi���� ��&8���db���p�唕�?~� =ǹ�����Z+/$�O}ȳOT�� yDvnI�Q�X���Yu
f�]���V�5^A5@�u�Β��-3Ù'��@� q�T��g";;� `���v��b��Uy�����.�H,7�ua�[�4��ұ�þ�$��ϋ�a`��P����j�q���[
=#�L��3YJ5Ⱦ(����o���{�x���}�Q��;�Z�K������/ġV�ΥБ���phMΞ�q4�ąTbk����ƛZ�M�� p� ���wOO�l|��ZM�B��!�%ڷ�=�Ll~���5 ��� ��3h߸�֗�h<� ����鹨Cj�t}/zf���̀t4#~���P�!UB�X��6	��K����=���&��,�v���-;�e	�r
��uF�e����`�|���o�O�����P�9�6�W�RI��Q_�m���C�:
�������2ٶ��Z�U��S��\SR��#<L�EJ��y�yM�蟹�}��M�{�4i�2�>�|V4��].�B�y˜[e����"t�q�_W|ȅ!u�U���8��Lmm%55)�_���������Q�D^ޟK��T!���8Y5�����@6����
=���g'�{W57��5U��vil|{��-����/~ �&��⁢Ǐ_��>��T=�����Z"����5��#��>���o�1�J�[Q���|7n��>N�_�	�f�]�Zm��� .�'�$`����!X�Q ���n��5���X�t�z4T?"�T���,��2$��K@g^������h
���X ���r����a�aLH�e��АÓ��p�r�8�rnccc�u$Z9��$�Ӕu؄7� vf``xY+����a��[?��ɇ�V��� `�$a��ڀ�{({�b�����UFɔ����І��Ng����������[)�p;"����ҷkg���|�slM���-�!�a]e��>>�@!��mU�^���0�+�Qs h`����X�J<��c�0�}�]^.@���tfSvi��j���/�Å�[7u�;�GB�WM^@ɿ��Z)8<�7�r�5��8�����,s5��ҷ��,���M�@����;�œt�:���Ҳ�����pN�tT&�}�~mt�(X?[������j�¤k��M���#����+�^~�F\i�]eGj���ߙ�,j�8�|ȍ �իW������d_(q��xω�@���F�~]�^L��������{MK���><-�&�4��4��K�苖٢QQ8���%�cOJ0C��g�12r58����텇��,�pa�o#��絛lJ"�n�>�tF� ����JS>��O�@�2Ny#=�׮#�!�y2eM~�(�,*(�x�?�uU+�=\�������Fȥ;8�{�ahO�'��痖,""�O��Q���'�T �E����h@�^����p5��H&�TV�q�r���\MG�y4w��V�R[�=�b��a�I����qC�U������lH���}�|!�뒂Z�t�6�Ԑ�U�_̢cZ� �����S;�n��.����j�CVҚ'"̊�1RHT�b��죄����Zs��س�I:�R�%U�%�E��섄���)p�;v���g�H��������2��Ѵ�Q��� ߛHUn����@|��(��6�C�Er�^/_uQ`C�7��Y&0p�_��p���P��*dR���u���!>�^������	��k�,�^yM0QΦ��RCbЩۉ:?��6g�Nܱ��򍃜��_�Ϭ���[�93lcE���%^����	�܊�S�ڗ���Ԓ��#-�dX.�j��ȡ8״M�Pj�{��� 9����YYZ:��t����5m���7�&B�B���ˠګ���y�ܚ���*~1�O���j�`*�F��Onz�,sZ
�%A9V�6�,�E�+~��#`�r�6a){�������^,���
(K���f�~���. \���,��ڼUUgۚW8O�z�?���X$�c�B7?~� >��e�5Q�驏yB��Df��I�<�KĎC^��.n�C[�U�xC���g��l�`϶����a��{k@t�	Fxxd��_��h���u�
v���rHc(��z��̣���4����Vm��E�մR�B�02�s
֣�߰��C�lWn�\�S���#H��s�{�>�M6(�B Y8�;�y�>e#�>}��l�(�v��	`�g�%1�y�Kp�T����<Û#'���A���a�!�7~M���o�zj`mt������+t�����X/̞�x��%_Dkjqkj=�y�IJ�Λ�+ŭ���u^�5Slp��mwww�����{�](��G�wG5�m_QP�*
*M�WA�tD)�"�z��Wi��@��Co�ti�w�Z���x�{���;#��:��{���<g��.�H��7���Ձ�'�㇛^G&v�G�z��mV�u���X�A�C>sraX$����f��"*Ɍ/@N�8+����3i�Z}� w�j����g�m����$��;�Ȋ�i�	���˂��l��:�y����0S5��ͅ�Ψx�D��-99y ���M/.5
&H+mDx���y �@^?J � H�p��٩��1�tM5�9�����>�/W\�0���t�ޣ���vu j����>��8$K���A�%�DtC=�&�>Ѡ�?ծ?d=�o��W<_	�P�5!� /����̄�����Q�A� ��ҶṺ�����k�U%L�=$�g1��؏>ܨu���M�}��@�y��
Xxtm#�s=�H�!���&~�r1��=mξ�)S�ֺ��H��a����/�dn*����x����GL6޲X&��ȪC�f��j6p�����FjD�ڜ'�t��S��JJ��O�`_i�kul���5\u&{u���Qo����1Rg�0mVO�� F�sO��6��WQ�jW�^c[(Y�6˱4!����̺�}���WkNM(�
^���<x� �q�$1`��@�;��d��8�.E��;[���t��7:��*��'��#vD+�XEE���u���o�ݲ]��H���'%x�:$�p�m�06��gYh�o����y�Ԫ��Ґ��(]�΄�.gܖ;������ׅ��zd����]�!�`hr2����}˒0X����cڠ>(����U������0������8����%%gr7'CT�� D�:�M`�n���B���W%>��SM�Z��"�[8����Ĭ�ri�ٴo�����^�a�}Խ�*лt�`ƕ���m.:S@��(>*�D!�/�\��ƻ��TB�oo\��^���/�*��Č�2��´_0�����#��&�rUm�r=�X�mOZ��.�a�G���:��Q��Z��獰����6��Q�d�鱩��:��&�Ǐ���WH�~�-�r�z��H�%�&g��5����Tݒ�����*��c����缐z܀Mn����r�@@xʗ�d��2<.r��9˱������mf�!�Ɂx��]��͈s�9�0�]1��"� d0aL�k
&���J��(�U�H `����K���g�� 0j��jmm��~9��t�]�~���a3~&0p�N���o#��P/��H|��4��O��tu�,G�X�����R�PC��i1��p��4"�3��$%�CC,��ׯ�]�s��������C���-�PC��Nn�#ڻ��%�Y��7�.�M��:A���sċ-�>}�/���T_�u���k"�C�<�g\o������ram��5��C�/����o�Ex�nkhh�|�:02�[:ܠ����uh1Wo�b��j�� ׬1bn� p�F �B)h.T�܉�xA�@@,aA?2�Nw�5�%���^�>N�`����8Ghh�j�� ��!�]`�(S�3S9���w�׏����fq�R"�)�:�_	##o?�ց��mYI�1��Lr���0ĬH����	+]��0���O�H�&�~���H��ӻ�}��y!�����@W�������ۿ�ۜk����ȑ����yyK�,�U�;�Z�2��/d�)�$#0���@�X��Je^lF�d���� ��z�.� p,-��D�����e����Y$�6 ހ��w'��A����ېSYY�05LE/����u�.��_�|�~�������0)�N2����RB�"���Xw1q�Sօ��=i��K�3O�JlQ�S��)��-셓���3Ņ2#�;�=@~�R�2��{�qVL}Οh�8��ɿlW���h\�5���["��=x���zl|�9%$56:��d�@�Y�	bl��� y�Z��1����>�[q�����~~���#U�+Z�K�:�:B���TI_���1��rRz� �d<,"�#��ҟ�8A���x� ��J��m�	�� ��k6�2V����D%6!�?p��8�����G4�-]1gC]q��0Pޠ���Kݵ�f-���0�a^2� ��5��v�H�
��Z�n���g�֎�)���/W�h�n#� A:�Q�7���p%wO��i�i��W�e�'��w	s������^#�������hL9`��W�>a�!%~n���_���N���'���k_�C� �P��[G{I������`OU���� ����0�W�*�v�Oy�m�.�.�����$�����A�փ���t�m��ʣ+Cx�%���H�M����Y;���Y{o��������?�����jJ-��U���M)�^��,�n����܄<��FH@��������|�Zr����?�����1�Cx\0l��[� ߸Tݯ�������U!����kxnz-�%V)'V5/�)k��;X�� �ѵ���~�Bj�h�5�F�D�'AE./[g��&�5��@ٍH���D��{N{��`�����"Z�Z�i���h>��	��ar��������f�Cg��Cɉ4�r6D�S.��������i�H�'�o��q�B�D���^����1=;��`,Zjb��(P1��Δ
��w���A�*�����)�i�}O!@mJj�uU�3�у ���O ]]�d�:ұ�~_��Q��Чť%!�#)o�hE�ħ���M�D*�M)����o�~�z��y�P7ˮ�a-�ccЕ����P:|u�B�/~'��|��ˉ.��a�6E�r��::��Smdr��N��ۻ$��?b\p���Kx�LY���H��}Eհ��gFq��9�t�H�È�U��>�C�90�P�&���ob�`�cE�����r������4S�����c�*���l������#�=�=���n]Ā�JO�<���h;b^K4��M��n���E�~�JK�;rr�[bd��Z�I*�:�@59s�iH04���#�_�?t
�����_E_9F��q^W�����ǫF=bcW�Фl��/(Z[/��Z?��Xf^��Dc�g�Z�l�ix��3��L97_^Y[R���٨h<�����SO=���C��[�~WG`��<����6K��tP%ǁ�ʻ�⦧���f)�:&�p�%�1'��� ���А@y�3( 4��1qj�~�\�6kP\�¼c�\���@^A���̃�B�x�I`XbI|Z1�ڴsaK�ƭ�#F�;�7� ���{�_�A�:zR�	�ql Sn��+[�%F��c)��,ĉ�"�I��ib�5�QHz@�^�����O����Ǹ�h��l�=�&�|#�#ZQm��a?�b���ǽ[���h����[f (t�2�P���`��Ʋ�:jH�6�-���?�T�/Xr�9:�51������ˤzڂ7-@���K�䮑,p���"ZP_1�5L~qt�v�~�`��A�ݘ�U0�bg��g��@��}(AQ6 �uz���x�ϩ�)�leK$��^.'��h������%��Ռ��1C	����X�	4����I�B�=�߯/tm�"���P6��wy�Y��բ�D��5H�JLLLZ�o���hUa���&�
��3���Đ�W�o�h�+�G����n��)-8���@��-��7T���y Y_h��w�{��~O�QdpB��S�+Y�آ^??���h6�p�D*]J ~�Do��CgѠM�8µ�����!�=��ߠ����f�x���e{�"$���צ�ѷ��S��r�_Lv"��%�+�7;�oh�m��t�xc�ֽo� ���� |�����@6�K*����hi��m<๧�?���^I�^�j�����v'Hfm���D����Nfff��(�/ο�@`-hN�_�N��F�(�&�/W��p^E1�pQVL>��DT�� R;O)�P�x��
A��'��BD D�O��g+�v��DFxu�"+�?EG���C�4~���BXa!�e*�C{�TU_���&^i,v}�8Bg�4"�U~�<�ژ�J}OKpWB�<&il�8�h8�ڮȚ��jNd�������U�~��1E�3a&$F�"᪭���19�"M�3��	3���+.��ц���옗v	�c3�*<��U�����{���#�jL��%�%�C6�����6��j��+D�2a�}T#-�]-dj1M����Y|�����!�zkfڄlҩ�����bNB����Iָ.��Z��ۮ��<����d�]�1�/��ȯn�C����6���kʋ��|�\RNlQ>�H��W���0�B$����8I�O�w=:�!C���S��#0�j����w<!vހ/��ob/zxgb6��<��L4=a0;�8��|뢙�7h�ǖv�þ~��sO,*_�l`�ZiMI>C�^V<Zb�HI	�{J���uR�o��� lJ��bTN��������C��YZB
/��'L��o��� (K�1Q����'|FE)�|38l8PHj|x�8$.Ņ1~�H�#��x_��o��7����n?�oS�����_�����4,ͼ�&'5mC��j��I�ג��8k��C
 �4�K�I�+*�Q@b�͑�<�%���0JlS6�/~#�g`׵ ($$Cm�]/������aC�,���\zt�(�>*5�
>��|P�H� }?�A4F�;,S��T�p��շ��r̵����U��ۉ��n��dg?���K��@F<i�'	cdt��q2 ���H8Q�K�lF��~���Z�A�a����[��<���lZ�՟*�;]�;���
���̩��+:��ɮ�)������h�/R�?���po<T6H��܎j+�Sb9D��p�z �r\� <$F.�C90��f��}�A*�G�Y��ܘx�H�V�8%o#u��~I��ΗeiQ$L>˳�L�<����")U�ٹol��D � >�~+�;���2�\ ��܄��7x.3�sF�@�6'����Ջ�'�een���Q�ɩ���Lo�*#���C��a�ÍZ��M�!��+����<��D�֣� Ji���|�x�]г����Ӵ����GF\ٮ��g�7Գ\/������Ѧ�<�ĕ,�T
�7
2�+���j���r�!?����A�a�Ļ��Ff��!]�y[$�_@Uv���󒏄W��dhi-^ B�Е�j�X�����p���˲�ϩV(g�{��r�������ld���p3�l�C��R3�h�&�5���u�L���K��Z�Y�w����k�$D���F:���1R��-W ��tFCC�]�7Q��: [�]��^�])?�߀<6>ؕ4[��R��:`D��� �w��}r��T�g�)�{9�6tB�M�9���b�!Կc��<G����@7��*<��\0��9��u�P�?v)�;p*`M|���+������4P��'�����O��6A�7A����<& ��l /�PSg���:͋q��T"f�dvZ�7�^<�f�B�}��N�h��-���&W@Bn���,?<G�T����f���N�i<ف7��%t�o�n)c��G�aVYW�P#:�j<	]Jy��F�Z=� �M��� ���ݨ1Q�`0�1�i��"\\*ܙIR���M�^�HJI$(B�f¨����"�)�S����E�O� ���8�բ
q��  ��t�ˊ��;b��G f����	���2
�O�`�X�s3тt�r2�.�֢G�ՏZ66@UVMU��%��\-�+���&,��![�b�vll��k�r��25���:{�芥�Bv�y��w ��M�y����^�]���4@}���#/��d vO�Ӑmྲྀ7����nnn���^?�g��d7 �����������7��s1�B}b��Ș���i6LB
j�C�� ��1�f��")�F�9T���1ZG�K�ٝ�b�t��������H}��cz��
{�d��f�{�%Ȇ���,�%����ᅊ>���.��� �ʹ,Ɵ�{��f!9O��]����pD\~1�#�q�hG�� ���>)1X�p� =�C�3����L].2�d�b����{�+�w ��m�"��/3��Q�������p���"�n�{�Q��w�s]�����DK/�Fb��B����)�b�p~�W�ϳ?��=.�����$r)�3p���q0ρ��H�O���.��lDmy���1}�)7B6D�R^�=7�G��s ƫH�&i�&x�0���Jv���y��[���E���2mT�F�i������gpY7���Y�C3=U�3��|3�%&:�v�ڪ'�7�STڑPi��ũ� �d~�-�=��[D/� �n�-���:��ބG!�\~��
���#��w���堁<ؗx�sa �-⓳�&q�X[ԭwI���@Ä���ld1�� !���dr4.�ԏiD[ ��)��g�Si_<=ۈ~��i�Zb�q�Ч��I���B<o��9�4d�Ү<%�M4Oi}���̞L1���ڑ�"���R�K�W�}\�yt����c���'Rw�t��<�Ҷ�M���zr��SSW��@Lj�8Y(֝����)���o�N�>��s��BH=˩-�o�L6$�+w߯�獴��٩�$j�~�!c��2��`���?��V�0�*"�'��� ��<s��U%�2��b�2
�AZ�Ԛ9�]2��eh+Y��f��)P�UZ������HHS��Vcv��8���� Oz�J�)��h�����-=ν�����nB.ń	����\�@=ٯQX����!��eL�iJp��;M�$$$�猛
���d� ��oȭ�^�h9>Wf�ۡl����L5�ݏG�)�25#�q�C�6��+��f#u��-�K?�(i��(���گǹ�Y?7O�q?���~�L�x��aw�	��dc�?@a0��C7VSs�F!�w1�����Zm%IH1k7���k��♏L[�؞\o{�Ԧ�Sџ��(�~���ȟ#:o���Xʭɛ�FO"��ҥK�?�0z��}\Q�����-�U!�����+?O����O�#f�9�Nȩ�"�pYcK�)p��c"��q�G	��tP8+++%w��p���s����@�X[[+5\��z9���*z��P6c�;-OPE���9�N�����d��H����>�����˝\Eu������ +��1�6�멹D7�O�@�BM߻�"�U��}����=g�/�ꛨII��gAg�s�h��ʼ��X�([ *��ny����f�U��Ǽ/�r+���2��_��2{n��!�=!��3�.��31{U�����sz�����'�����2\����$Mv���M��$��-�ꀿ��-�|F���D�)��V��X&��A��?�0K>B+0KrcH�=.����oX�B�ܟf���:�E�����1j��'�<uD:�^���P	�+��.����G�?񳶠R�A�րD
&�6�a�>]���Gd<iry��U2�ʻ��u}A}�fȵV��!׆so�@T|���n|]��)���lFkk�Q�����B��
E�ǫ��w�g������R=ryt�����ޱ� �I��ы�ܧ�C]�0�5n��:�f݊Y���mǾ��}ll4��- ��{9��ѓ��Ӗ�F�u�`���d��1 6d��
� �ۄӼ���g����e7��Rm74�F�.A��&p�U$�9����g-x�(�w&���N�E����`�TG{������x_��"���p0��]���G�r�D�ݵ�p�>y���A�om���s�N�[ԊX'\i�\?rTS�կv�2H@�X��.�f���k�����#�l�3������^
%	���E�����>�D��Sr�F��g��� ,����(��������O�"K�A�ӵ�V@�>Cں���?�-��Q�'!;��@���#��5:hM��	�}��g��,'Jd~��c�������_
tC&�.'�)���	�����e33JJ�G�㍏�_r��;��p�]c�?e{m3 JS �p����D���J� a��@�_3F֢��6v�6��������Ϝ >%桫�U�xKe�#G�V;ٯ�b�I<k�D7}qz��q��sj%���������X�+W�dH޻��Μ{� hɍ^��0�R�1[U�ͧ��q�P���'���b`��3>g͂�z�oɓx{�E}}�Ҁ�;}�[�.j9��}�km����w�f���&6�����V's�G]�xP��D���<\��o;U��]��!9����Lv��v����[e�+�o4���}�!�S�\��lE����g(�d
6%�?~,��+C)���'��-��󵩮��]Ko3�A���S��DT��Q������bѦ�"2�	wO��ē��a,���3a�#f�)J9���&�����A�f��΅�ׯ_�?'X"�bxB�K���y�Z�7PnK��5����+s1Y��X]���{)`�<^'0�qp/��_0r����=�(�V���ݟ�i��q=���7(I��c����pw-ޠ3�k�v����>~� s�d�BNT�K���4�{=#�3E���TWdP�)^�w��w[�C��K��X���I|�;�Aҭ@O�X~��vݿ��r���s�6bR�]�a��F���:�#&X�'����qG�RXҬ#Rr1��Q���(he�));i�5��q�kޖ�R���h����[A�]���� ~jqڸ���Z|5#�[?T�HO3w*�l�V��6By���3�)o:[BW�om俼ə�܄�	�U&�j%J��.�bTg��un���R2�=��۷oY���l:��[R�Eﮍ=�ä�u���96!�}��(��}q^����{�k�{ON��b,�&-wl���7���e����{���y��D*��x����M���V�լ�F�5H�Q(�����"�V�����T3�"[!)W�ZZ���K�G�D���@��~�B�n��T6��CRR���p�ѡ(����(|���/pa^��0e���mxEo4�H��j������Y���+g�ҼId������Q�����,��W���9S�,��-��g�3�T��J�)��*]}����!Apq�s����Ϳ�c���Z�|)�|i�(����&:�s�,��²�7J=��eW���ݎ����}��߱W�6�����A �&h�6����X�!*<l��.�'�S>���rc��܏�lB��IO�=����D����a<�z@������ӑ��&�H+@�ThӇ���[&�RD�8J}$YG�<Оy~������=��J��/��qy�q���J���6]}#�u1�|�$�T���	5�'&ބ�`<ˊ��Mx���ڜ�G�!�T	,�����O$���7�1hΐ�_��T��*=a9���+x�� �2vȈ~����Z�Rut�8��B���E������'��}lP�N懺S��G�؎pL�;�u�Ol|�����A��7���v	hh��(]��c`�	6$����9���%NjrU7���B^��7OU~��qN�'hOftƀ�̪>����]h�N�;�6���F<�e�rf��*���0ʌfh)�w�R\�¢RH�$�q.�Qʸ!-'�|z{(��3���6A���F��'��Oz���z)5���K � '�YJ-��;8\U$`�?��Ml����ZR�K�<}D MN�i(lxX�`S�y��`�`̀���Qu;�f�i<��Z�H������~7"<|r���]�3�E#�}TK�`��[��⁷pt��4�b��i�H��.q�����(Qڥ�0 ��r��1��C�����:Gf�'������S����R��O13e�/Hf�����+��/u�G�%8��xυ27f�@�tmrU�7{Xh!��0�,T������<��Vǅ�����Ȏ\(�zC���`e�y�O|���V�矶)ڲ3ߵ�k�Kwؾ`T�/�#��H��}�3����� �F�0x�>�:Ǚ�u}x�G-nM�Y�8G���c���|@�D#�In�/�zT/�*�R�DW��:'�_9�fڗ"d{?�n�S��tݟ�-=�R��������J����(T�aL�q<��r�� ��`*.�b��(F�-Ne�������Z�~������)���T���_&��i]�ϔ]��t� ���]�(
�����Ng�S��<f�Ԗˉ��o�̊�<�����T���rd������>���|��4ہ)l,�1T:��P2d�Lp�}8̧���'�)��Dm����`a�m�s=?N`;��V?��tCSE`=��K��2��Z�-\/�`�GZZX��U�{��%4���Mx75���G���eB��_���a�Ӎ"*ė�,�MR9�{�=�ɇ�_�f�����=��� ��p�?�s䨇}���׬�\��Q]Bm���A���J�W�c	�(��p��wa�Ú�8�-�L�bצC��W�\^�
ag�ߋ]���ͽ�D\�[��{���#���o�ǩC����7�8�tN��k*k/ m�d�H��dPs�*mH�B�H�6�χ�߯�uK�=��Xiz[��c-�6-���o�O���n�G�E����Pl���؅ �f���c��<|/��Ҥ�=��&;��͆����yl<j�뽵�������۵3���{B�03#���3��h�rhĵ=HA��f��)n�޻���b�uo2._���n>�_�5H�QW��C4v՚�8U�wQ/�9EΫA�_2Gsd��~l�_a V}%���8���#w����@t3�^��7�]%�5;�H^�b��3����'�y`~>s�l��FF���#�HǑ'F���p;��5c��o*�1Psˊ|� ͅ� �+c��'�@EtØ%�n��Y_�ڭ�Eaa�R!]��Y72�/ad��aέֺI��1��T�����o��^�i���x�%BY�s4��b�*�q�*$��A����jQ�|�;����'�0V~�!:��s�����)4Y��հ�6�Kgv5��_����c2N�WW�c���S7�d���}񹔆��\M��*�I�Zq�w8%�=&iߧ�?�&�w`��R�e���XA�|Sx������|�]c]o|��/�.��ϜP��ߢП�gԌ��~�m�=��߶�R��]���ӟ���"��x�:��|<����'iy�(48������]��������7��&����
�AbUX1��Y`�=���!�^3�v]�SB�?bD(�&a(�uf!���Vc�+j��a3�H5���U	P��l�p��7�'���|VXHڃc._ׄT��_;y��	��[�%�c-
�}Hۈ	�/HwN%d%�N���0�q�`�y��NK%�e��v����N���<{�����#2q�?�-Fsb@U��(�#�@����}���l����ۜ�n�O�	x*���%yfk�֬�Z���Ϩ�� �*78�Îb�<Z��i_Ȩ��h������k���8�Fq��3`��=Y���p�����R0��갚�ḃy
�ˌ�]W�UT��'!�F$�.��.�!D��U�9.��R�@ڗ����|��
�|����Ӽ��_�>��{_6�nk���j���	�����:A�1���N��_ nK��=����9y����F`;�^`��Ⴔ�B���L�o���՗�4�$�O�s@q�뒵���ꍂZ�%±�0���K) t��WY���R�F��'����������,�t�f�gL��}ڬ��6�6�Є�)��E��
��U�6�8WE�}���au�����y��fMě�l4����/ƙ���QZ??QD��, 
���]���{�L�q�����>?���4v9X�ɝ9������SK��+n�x�a
�d�嫯)�`�r��4�2����˶�ҙ�@R�J����:���������~Bk��(��<��洮����ɯq7�%�vR	�3K4E�c��N��؃�<�U�!�=��M�/���U>9��w���:�|_瑟Y�J�y��l��pw�x���ȓw�M��&�q�~�k�B�����Z�^�m�T�3K�*2H���Z��N�9��u�;a0YN���8���s�s��¢n��J�ez4>}�q��ٿ9*N�xP���*��s�{wAe�byܾt��w��r�bk;m�G����wZ����/���Ο��R�_8x�V��V�q��Z|�N�K���=U�����/�S�oWEF�'"�X������̞Lw��|*ӥ)u�/2+Fq�ǫ!��}�ǽ�z�]�c��AU˺qK����ɒ��3ݱ��нR�u�}�π�7/���]���d�mՁq�c��-��=k��J�٫�5h� ���Y��r$TM+헿ךlƨ��=:����=U�"�n��Pem�p�
1B~�x#��Ke29齙�'��~�H,�V�Ԉ�m�D�	��e�_���Q��5��)�%���;�0�� (��d+����줯�K4E�0��S)�Ǜ���Sw��h����PoI�v��2��#{oI�ԫ���*�;����mh,'�;�S�n�F���lM����՝�ӖC�pVpPj}/Ų���$|a��(}C/'B�؈��OH�jﺾJ������G=0�3��Q��$�zz�]��,nN���R��f�Og������DLC�a��A�ԓ��̡�aȡ��&]����C�� R�����}^��#�����Vg��~Tw��W__K�V�`'�?�>�*r�%���n�M<���p[$��w2?`�7E�zb��`�|�������5P�	��l���bu׷A9���/�$�?cʡ�u�^(~%m-o��6��������%Ѫ�8F$p��*$�|18)h�_�g�Jav��C�Vi~J.vR��7f*_�G�su��ڻ`����s��/��
�|1���*���Q���@�k�T؍��TW�p�W��g����?mP>�`z�y�Gڐ@B�_巣`4���Qۃ�Z�;�-:�1/z1��p�S����JPK%�$�!�������������>���M�W �F߸�����ӡYS���%���":7]�~���>�f찥��3D,����ٰ,p�,@s��`��_/�Vc��%����U��a���Bs��Էa�r�d�c��絭�#�F��L�ۧ��G�2F���
-� u�}a��<�P|g,|AH�!�Ɣij���6��ĉ��V$��]��<6�.7 *��N>��k[�c5,"�u�n`��<5�!5�o�����<d���z�R����P|��8�Ɲ�0���N��$��Q>��z�&.�o/߈�Rئ�'�d,�u�>H+���бƮ$�����^>cC�m̔k��p������U-�,x�L��b��q���o�A?g�������юh���,=3�'`��<��O�ϝ+E��J�,�+[{|�������V��xNF����Gm@����`u�X��o�)�m�����&�P_�,���`�9/C�=�g|ݸN^C�������*�-9.,9$��,������W��OE0Vc��n��k��4 �ԓ/��	&��X,�W�*�r���뻗8�oYG랉A��UBB��V-�#����˜��S_Ɠ��oS�)AH'���Ig�b���O�������`�l���;r�7Ի�:����m�m�:V�jQ@"�ٌ���j��UJ?>n<\Q�wy�X9�|�&��)4�!��2!mw����fO�G��}�����UC��Coķh��Q�mhj���[��s��)`��N�tӗż� �s��OFE�9p�:(�������l_{=�F�?{���_�<�s=s����j��&���R,�#��s��6�ثAM�FEk���"(��*p�p�1��~0�7+d\a���u���������p���*kڂ(5��m��J�3�#"~��?~o�k���ŹXP�Kŀ�Vc���V�fm@���'���Մ�u�@LK��R>�XԻ<*�$Zm��pX�5T��ߢ'm��y��w�B�1�k��²��⓲�ǯE$DN�f���7K
˸���{[/���6�ɝ�����om5��6tⵌ�Dm��*'�K�ޮ���jA�0�P�Ju7�,��;Nq����P�a7,��ȖA�Oٻ�啘�i�32.�����;z��E1U���]X	��������0~7u��N��2�*��{���A1�?o7d���z������v�/�;�h+���-DՌ�"�ޡ�\IG�Ϙ�)�O�j�U7<�j��@K�R!������T'�R�-�������X%�D��][�����ӭX�T4��Y�/�M误u䏓Q�>o^�U��X��vS��h��~���I�`Rt�w�g�͈���Y�����/#�3ƿ��wMx�1Z�����nCF�U�9p	k�=���Zc�Qܺ���ZtR��v�:}Cl��d��4��^_]�Ή����D��2��?s*���֭�Q��9{;l(R��Y�����#L~��P�\��1���%}���c��+�c;:	����/�vm�<d|vC�(O�8�t��˪�&���!���(��B���>�"���;$8흩X��Ŕh�缉޳�C�;�Y�g�p�D���G��V�������O�uy嘘�:,i�׼�䓊�bAz��6�ڿ;84����6�=�*��D>~�c��d&��p�.��P��a���r�U�!~�eͫOi���5Kb������CY0P+�[I��B������_=�U���*i��o�|�pV$���º�L�b5)�Z8Q�4�Vu�z�f�8]u�*�q\JP��J�*�}�0�\K�O0�~��P�����O �qY����o�W+��i_�ܜ���:{ ��mүуL�P�Tx�>�]�0�s�Uf�P9��;�����=��SS�|����r�Λ_�&����&�۞�]�]�l���,�z��C��ɒ��� �͐g��C[_����X��{�J���k��rwN�&�6ė	*��n��A"J�Z#��os7���jy���\�t�:�c��_d���U�-���Qo��fjLP����U�XA4+[�q�Y��b~�����qa��'2h�Ġ�ܻg�e���lY=EA�2����F-{�lZ��l���������w�_R�1�3��>%!�6SE�"��ƹ1���ua�>�xːü�_�3�-;��s%4w͑��1������P�n�}�CJ#~�1���R�E�;�>5Ξ�n}��q��"eK˄�eF�͛�Q~���bU�^���/�:ho�u�p|�w��zk�E���q�a'qO���ɬIcnQ?����"��q]3��R�)l�U�׈%�hD�����V��L�z5�ŧ� ����WC�pZN�gN�М�g���R��ɭ(Y��ΗP�_Z\%.�|"ehV�ST�t8׭��5���~��\��GI�����:�_���Lk'�-�LP>z\ɖ�9ob�D`��/ף2�T��9�:�h�=��ـp���e�z�n������h�T�G��T6�q�̞HY@���jo\���}�����Cv��d�x�.�d%1��S/OK54�$�����G��3�\����.x��y��ͽA�Y��w ��ֲ��US.�D��s�f�?���X�;=����o�0��	��׈&��F�����N�T����@�2�NRt����͡����/)��9s�
��&��Q�u�ǽ��(��l�8��t|��k7��������]��_���ؚɂ%�b/�z?�x���5�'9ƞ��w�N��6n֬;�FZ�Dd��\,�)���ʠeP�O�����^%��SCbڜZ�`m~���r\Q�(.��l`�b�91�8���P<$%q*fz����G���>��QB�*D^q,�M��<�$~���ɇ��R�D&��t_�ת l�2�����mQT)ۅ�u�K�e`AUtQ��б�χ�M���wR<}������u�tZ�[+��
��s�JJ��D"�r�?�0s��{�>^�/���|���,^��(�{y�?���F�H�M������I!���������\�i�h����*��;����N���(Rk�'��a��_��0ń�Ft��t|�8��gz�V)����(�aa^3��mt�L�����]��B��U?1�-���#��%�PoY}�{��6�cOQ�/�41�f�Ǧ�ecg��l�>2j�Z;i?��WqǓx���'ٵL<� �U�e+�1J�K�T���R�;D�Ƞ)-��wF�Z+U\,eMd֏4�_8MV�)o��o�m��� |��!2��ߒ)C;eP�®�k�[m,�T�)3�V�6�?>�y6�3vA���;���܅�ѥ��*�8�^�5V���{�;��K�	zП�n��u��y025���/V6HvƿQYu�����C弟�`N����1K������,I<9���|�z�����w�a�(1�ŭ���vy�d����]o�'R�`�k]X%V��%�JQgn	�#��U����N�l�����ܢ�ء�<�JfE����,��L��"�h�EW��@���9�pNe�.Z�j65�ٖ����:�I�R�����b�ȱ�����[���O�ڤ��y�L���E�~���,�h�N�N���PR�{��Ĉ�`������Y���7��qUV��{w
b~jr�
���u��-�i�:�9d�.)��+����eۈNt���Vqvtnw��V�3F�u�=m`N���Z#��|�7\�[��`�X>͇yWMl��0V�9l����t�M�g�r��ʨ��O���0'�)W�j��v��\��M���V�/�(��<ȃ$M�Мq�ʥr�%�U'�s@�%��ѣ݀�elˏn��,9.V7�z�S~L*��O�_ �N׌vo^+5Aw1�k���#yS���wh6���	�9_�ԕ\�u�$��o 7��I5���GQ����+ 9�QrO��ڟ	hH�}��/��\��x��2o�� ��i	��j?d�u���X��%!ɚ��c�p���>s���En�0��$8N�=�M��k�[��T��>�쥈��×
��m]�)~�H��ȑ�~�b1O��:˱�����>X��8����������lf ���{ϰ(� \E�EPTT�
"�!LdQ���$�!��dA@�"   9*I�HF���3[���{���{w/�9g`���ꪷު���\&�ڦ��������~��˹��
�'���W8�O�RE�ei�tI�ı��]��g��ʝ��^e�g)ݫr��+��gq�d��%@�C-����5���n:�|�+W�MC�BSV~hI��+6B��@���%���A��Ky�'�+||��~ϟ�^�ksJd�d{z�D%z{�'O����[�-y/L'Vx��2�P�-�y�}��,Ǵߵ���6�4H5Tb���L�$ne���b�Z$�{3R+I!�z�����'�m��UV������ Ý���u��S3�nʞܬGq��Z5�M܏U�5����%��W|�`�v��<n�����薈k���}_��W�3S��<P6����d�VVi� ���m��.��=����h,�����S��W�B�OP;�`lmCU����뫻W�i���lJM�5�уC�ɿ5�y��gR3|�����+�f�����3\[�?ݳ�=r�}���������']/)���[�fh���Ҩ�M���SO���[��h�W��� ���a%٥lǕKvo�V�P}|������k��n<2�U��S?W��s�����V����'Nd�o> ��(��[g��K�9�L_�2���-H$���S�e��i�J�9nm��F���<��%�W^��\���\z֢z��}�=�IA�{雗��!��
�6����Q�z(7��5Z2\�bR���M����w���X��	�Hާr>��+c�ƭ��L >t��FM�`�E��^�k���_G���J��zs�rd �7��-�Z�Oj�4[�<�yJ�����V�Xu�n��m��ʢ��ql�-"����FW����7�טZ�,�5�,�FƖ���g(��nm�z��=9*}C��<��'�i��mO���di�Bj�q,%т9o	��v��_}�"�JhD}`�_��t0�|S�"[��&� �>�+��W�S歼�C�s��2ç=���q��h�+;!�m�����r�����I6�����X��Ӣ�OE���|`����͂ڝ�RKL3$���O�
��Szn�ޓ!�ם"��[�[S~O��%H�ɋc��'�N
_�M��Y�t�|U~N�]�߉j��;3Gy�;�Rۑ�� [�K�7�6�A�%eu?���h	���^n�:'�5���#�3��+j�4x�F���GG ń��+�5�O8.���������k�o��D2�{�E|g���{wi���,4~����y ��� ��:��/χ L7\�7����J���3|K�D�5ǹ�Ж�gT|�z���x��hZy^�0�Ǚ�u�=��o��~�n@p�͎fhd�j�56�h}�r(���7��}�fRʂ�Ck��e~o�++,}o���vxqP;��U�����ǹgߙ�O,׷����������N�;V%:n����8�asنr׾0���ë�[vd8�����.vd��u�E�K���1y��RH��.�ĩ���*��7<si������wr�I0��ZQ�ڼ���Ϲq���� ��[�4:�}N�[/z/��s�Ӊ�It�dN�*�n/�̻0�f�{O�]ɍ�����
��D��-[6f�F��2��?�>V��'��NX��$�(s�ߥLz�=l�<�6f��#~׾/����zG<|4b�\=�E
]��Ќ���<|�b����Sz������a�ƽ��_9�}����bQ�ѦS7�͟�S�h�;e7I��v��;�O���^J����o�K���͙'�]X��+���?���S.�����H�:�w%��;4J8Q�?y�|���ע�!�&X�Lh�o[!?P�lq�C�Oݏӹ�'�D�}J�9=��</}e���w���}O�};rY�e]�3��l0��Q����}�ޘךϔ�KZkr���Nq2�_z�p,�߲���,�������	'�H��>�]s}��9��[����W��W��On��sU�n&m�������:�g�K.�,VtF{�*01�-Ŝ^C�Z�ރ��5�oH���O�V��t�|�ؒ�woU�>�c��?]J&�=��d��|q�pCV��v������_�z�L�U����l7��&�]�!%ٝ~_�������+�ϾԴ[5�mE5`���뗛��ľo?�m��Ή�į�*?����۱:xF�髯��"����Jc�e���ON�#�������}ږMۙ<n�\:yl#��MΒ�y�?]�,f�1��ʱ͗_��sYS��_1��s�(�۶���fP�N~�4L5��V]�RH,�7,<�����F�&���I��w���AJ�geVӺ:�퇍i½F
�%
Dw$�7��(��c�"M�;�%
��sVT�Z,pqCyKsó�;�N�J�Q�
��J&1�<m�*QN����#�t�~Z������[ڛl��Ժ�R��9���3�c�����LVsg���5�=V���:h|"��zL<I�?X7H�~JpLs�̴\hg>4d�h��3Y����K	��{(a�E���M�6�#��b��	�ܶ��_�����J��H�*�����[2�.�ʝZ�d\�M��,�pƑr,����ˮ�+#�������{��������]|���A@E�5�F�hOE�81qo�b,�.>�k4�G9f��{�ݗC�
��R�:��D��S�i�GJ�56m9�1E�x�tT������7SRJ�x9��hIF����S'f����9T����b|�j�S������ܙ�./�/���O�s?8á��c�N��n͍r?����~����S"@a��]���ゃ��*�^`6���
�S�5\���F�sg�<�l�ݶ�j��
5)s�ۖ�z>��d��n�8��c��@���޸����.�d�"��9�C9��?��fi����J�Y8�{�&�J����9	�iŜ���#�&�<-�8���^����,��Plq�>�lyZ�~�H��Z�-�cm�6+�3�q�z1er��Q�Q�������D���T��kdJ�vf�>X��<�T/T)6\ju	��d*&���L9�;�30��ޮf�MC���mU]Z�!�J��}�-������Z��à�Z'�A�e��n�!1N�)�������� /L�9{�!!�^��3l�Y���.'ǩji��2�ތ��v����X�<�9�:��n����Ie7)�����Ws6H(�f����MY�Vs�¸���a�3�}�G���˴^�t�՚�/w����۟�2�,�qϲޜ�&�����|E��vYtC�n˔�)A��M-�-�5����H���]��`�i)~Gmqt7���;��2y��Ȼ�ߕe�Q�dO�u�p�гTt7����	�B�吗�����К������6*4&
W0u̴j��|籤��(I*u���>Q���+vw�^�u�mlc6�� �M�F)�������em݆��w�#��i�M�F��H��U����e�����FB~	^�����NL���j-�`Z����c���c&���6$��3L�LԪ���h/;LFv��z�}9}���g����$z7�*�פ���
�+��O������7�?�4r@�5e��m��N˦a2���]�?M���1�'�u@J���8Q#x�;[�}~�5�V뇅���WW��R����$u�:yTװ°yOot��^��-hL�<�n��M�Gh*��d��-n�[�Qy�o����>
�b0�ْ+4�B���@q.p�e�g�=����[�lI:����c��;9�i�bI�N;�l���������P�tQ4҃i��$oF��_'��~�uS�}���`&���Mf(��{;���P���gϲ߾��}�t��g�6?\X�L%=%Vkx�e��Ȝb2��r$W�s�G?H�ّ�2��W��'M��i`y����!�o?��3"��?������$��Ӣ"�5�R��]Ф��]-�nl�J=�k��̍�M��d3�:[�4�<�����Б$�7_���������<cf��V܆��P��3���C7Zw5��j�(`�f�d#�N�0{�Շ��֎�*��\��%�J�zu�GD�TFp2�Ns�VG\ԃ��־�c,e�������^�`������6�Qy��u	�_��Qޫ ����{��y�"y��*S�p	Ec��g����7������(�?!�yg�-�����ݯ�����+ct3[H-�Nw�>����^Pʗ��H\"MńgK3zn#<g��$�#��ډ�훇�=��2�6�����!\o��f����*+�����;]/^p�1L���53:���4Ϛ�:MZX�$�D�����	�C5�	�Ő�6�)I�_�A�~��&�~������;Z������I�؃j,#�:D����saN�V:9����ī��J��_�d�|Wj�2�>��mԈ�E]�~5�g��J�ͭ� E���j�ڷ��Bݐ�V�@�|�u�P�nv�k4�:H�)U��G�)�vɐ}��L�M��k�!)8�����st�;Ty����=)�3� �Q/�'V��^���gk��q�B�L����P������|�iG6l��oQZ&�~a����{����w��3Z��;��fw*�i�Kp�Շ�˯��ߋEI_����M��F-�]�v�)�mF*�Z���.�0�T����g��E;�?j���|cMgǴ�ˡ_�5��>E������o��Ye�33�H??���l�i��5�xp �)����?_�F��g*�g��rMp�;�Ln�d�2�MQ��z�&��|��Z8��ģ��ޟ���	;�w����ۆ|`�ܞ�J�d����E�]�_��N��o�������]^�.�O��'h�z��X��u��"�E��\�.r]��U�+Uq���|�xjP�g��G�{~�����O��?�Z���i�����O��?�Z���i�����_rjLL���Y8�q�s{���[g�Pܣ,xGⱑ��wS��iՅ�މ��ֺqqI&{k*=��:��w��S��������T����x�ߒ��~����,��������u����\�.p]��u������U�G�	�#�b��ȓ>~��ӄ�F���1S6	�o�"�����y�>��t?��(&�md��]����2�8,���L4,Mx��Г�ݽ83S��}Bȫ��S�P�|7�͓��V�D�i�H�Ȭ�Z�xTEO��e��,6MU6J����2U�`J��l��ϯ�eU�.p]��,0�?��]6��5��3��RV�%�Wv�;,�\�������̛%�/�g�_�5�1]֤>�g��1�ǉy�B�sU��|��ݨ��v�8���#}�������Y�����br����ݪ|�̌q��k\�.r]��u��"�E��\�.r]��u��"������ �o��gb���Lmm����Jm]�%{������a[��Xm}}����B�b��*�鮮����\	�� .��� .JJ���>~�~�7B�g���.Z�k^����7 i�E�8w�N�g��[{<<<�~~�/�����+./_3�0??��cPa���Ϙ�(� TTT���虐�p��A75����t0��9�����c�߬�����ի��������ׯ���	��(��������S��TWW��:p��0Hx1x0Ix|~��k�g��h��ٟ�;��6 ����64�c�>��~JN�dkk�)�>~M}�%�RU�16߫�||fff�x|���,�4)O/hβ�A�@����`{��A�F�mҮ`�dɻ���X��U����xCMMm�×l��zz.h13m�LG;[��LgG6fZ����[�.�|����Naئ.�677���:WVV����4J;r��\uһ�����V77�y	�_s��(l˶�
4�qiʹ,N�(ަJz������6G+�%�oJDC��i�_�	���6h�52���mc�\�|�zC�J���0�Iǹ78˸^�ձ�E�8�=�N�Ŵ�P�z�ko_�K�Y�~a=q߫����9Ϝ�S���f$l�^$��*���F2���;������LNM]266V6-�wI��XwE ���Ru{;�NU���쯗ҝ1�9��˳�֤�������bѠ��jN��ąߎ�/�"*{3<3���ٕ���Ƒ3{Tda0�1�XVJ-LzI��A��(4K�o%iK~������c��Yk�E�Qk2Zi�%n�p����%i��;���'t�PʹZ�M��W�+Oҳ{�f�:]�;Ǌ�T2�[���������E�|we7ڣ3]����08����}�+�|�����HfOz��8�aw/�ypL�I���;���8�v��0r�`�綱�Wf�~v�|(������ܯ�cs=���C?��O��_}xT{X/V.J,Vh�Q���Mu�~�Myy*��8p�?5�;�F#�+9�����9b0V#����{R���J��A�R����;ev	d�SS����`w�s�����
ܙ�ƽ�lmm����000�6��Ps�I�#��->w9��ʪ�3���B�.IKKM��'��}�9���Z���M���y(�Z�uHPa�����M��1�XĦ}�&�)5�F��^�����lPs�<����N�3u���D�#�@�g�/^����l�cӕ���_/���r���$�R�ӥ��m��$iW�N4���S�u�x��2�\!

���ݢ�q$u�)_��:|����:Щ��S��[�8Um��hU��
�ۼ{�K��D�U�@��/O����XJ-��9x������0�Ϋ���p�̞is�M�/�Y}z�����@~~�i�$�>aR�y�����:E�C�<�B+����-a=y�5�>� >���f̥*x�aa/B�ͷ���vGQ�F� r�h����;�[Y�e�������9@R��?������W�up�r��������E���B�-����Ѐ��{��"�6�܌A��3��%�%��m�l��K�Sc݁�E<����09M�c�8�T'I��{�޹P����~j�����n�t��]O�I)��;�S��F�!ŹRX5���l��v�v{�j���6��h> ����۪h��w���?^WSCe�=u��0��mߩ�.��.Dʫy')+/3������a�f�,((�D��(L/W�cojty�]����׵�/f���$�L��E�~��m׽`Gr��gQ�܌e�ٶ薍ۙ�xf"�>�bͅ2��M�g�n*�,��aQ�U�/�� ��5ި�}/��\/��լ)�<��}%ZN�%JS���{�^-YY��'{����yfݞU"FE=�^%Peq�����~lz}f�UKz��U�I�<bo�J*I֔���i2�S���/w�ªu@Տ���^�����ʤ4���["(��d���0ĩ_�~���ɉ�*�;��<����[�@���U��l7;
_��C��i7d��v�1�֚�TΠM�)T�!�S[�o����H�L�n��lsC����vUH�fnN�Ѓ�O��M�T�����Ӹ�t_��J�����/؛��h��S��~�	KN��ne~��}�>U}�1��u��ϋ�/���ܯ�<�����:��-���E�~��=�2zʗ�Ҟ@���:��J&q͵��܁L%��k������A���wg��g�s��ͮ�Io��.�ğ�*��2�4����e#s���}r����eذ����.�P����GJ�7��I�
�lŷ�$��N�|H�d��@��[�K�DO
���:��{�awF��fy�WY�#2��^�mMK�b�>=h䬔���s.J���fө:E���Ϣ�T}1�3�m���O[��
��i�%�?��D����A)��1��]<��ͷr.������k
�݇��-���ݰY��~]<��(�L����8����Л�n=�[2 �w��st��9JcnaQ1�q��݁)� 0S	SR&X��!6&&�H�k�>}�$����tT�[�y������8�{�bǁ��+��x�F;f��r�U,nd�~��D�N����%D�_�CM�rvn̰0@�l�˫�JZ��Jh����� ��>UZ\jJJѷЋ��e9�Z���g�W�e��/]sS;��h�X!���������xR�COy�PP��|C�H��t�����奅�.���0؍~nL3�+�B����Tc������T ������_s���|M-���2u��v�3�ť�{����_׼�	s-+%v�/��+Y<h��8�c���pQ[�WL0�*�R<_{���tg½���+���v{qU�3U�F��gZ�4`B.O*F��8� S��������������0����{m��������� �3#UR���B��Ϯ| R��A� LT��J	�Ef���^�S�7i!R��2�a֨�▆{�5�ű[i&������3t+o�A%�7gy*��������N#>x��T����S ��Jݠl&ini�g�m�.Q�E�mA���75�:tȴ�`Y�'��;""�F-V�GV�ԁS�kW�������$��eO7ϖ*�xH!)�5�NO	��Τ���(A���3��n4�K3:=��[v@�ޔ���˪}���v5�bl�
�H`�≛q��v-Do���]�[��Ew�!�
r�����ٹ*G��ed]������N���u��ҿ�{�8�HU!$4~����X����%����o������
^�n2����:ؒΕ3�a\PH�F�,+x%.��N!~���*q�hk��X�,���9�KDx�xx�bX�g{�)���O����R@zh7b��v�#�Bc0"�x�|H`��m��I)m�:�A�e��:,��?M���N�x�������w�oލ�9����Y�,�3�M$��Un}x�G_��hG���EE��*-�u�}hT������b@�^J������q.��/Q�8��)���W{�oOň�瑟�A��񘋴X��}�<]Qg�[ס+	l���=>��ZG,���5#��k�E���<-5I��w�\��;s��M�ԇ��vghR⒳��Ei!5*�d}K�YE�.��*v6�WT����wZ�8M��vק��������J�����d����-�=q���~)k�~�m�ɛ���� X�|mꢽV!{��JA�7s�� c����e��vl= ɢ9~��]�N���(m�;�l��2�@>R�#5{Ȱ�vu�QZ@�sWv�%c�|��𸡶lfٖ9��u�MY�Bf+:_���z2ι���.2NŬ��Ӽ�� �M��I(
�D��.Ͽ��tu��Mo�l`�\�d��m�:�%=N�g�}u��+�\*�.�HIkf��Tٌ��7���yN�bQV����1���-������b�W��TLuM�K��_��;�+/�V����VU���J9I\���`fG��ҫ��4�fm��0<R�h��0�N\�BL�lc�H��(T{�]�i[񯒗0�w����|����"M�h��-�&ʹ�X-t:\�J$m��7��!t*C&;�w�}Vܮ�^R��O38��P���D5�'c �A��#������h-�ތ)�]��[xȲ��Gc�����%��<rC"�������ۗc�o��pRU��$�~yJm�'geiD'�~��P���!�6qo�򸼔���egl!�F� ��WIJ���Lt��b3�*����0��r|�u��`f ��`�9 *��w��)��4�R�� '�;
;��Y�"ӻ��R�"WE��g�۲��"`���T,[����K�<���Q��^��y���N���P�R@����=��J;��`�s��~a����{��Q�f��kF�����6\:��[�Nh��>9�����s��JP%��������^�u��寉!22�t���B�Q�M<	U-@<�
���|�e�㭳c]]����$y;&^���ug��� �q���s�A^M��V:ƹ��t������kz�y�v�;�9�^�u~��{,8����B���޾��+<���4@�$��`��.>��� ��Dۇ�� ��J5�~�WV^���*:?����]�\0�{i3؎*�M�Q�ɞ���f�7���X���o�%q�y0vW�SE�NI�>�cjEح\{<��00~�#�E�4�W��N!'[���Z�N$uQe������
�Ri7��^Q���/*�N@�8����Rǵ+��I�B��1��Z����dM�����J��������:��eI��d���,���{R��T��a�1*�%r��3��8z���/h��g���l�%�m��ݹQ��q�0�1�bL]�@#W�L�Vd�i�j��i����P&j��	��({���B!�Xz�=�~�m�U� .�"H��P������`,,1U4'h�}�D���v$�02XS'R��a�\����91'Ǘ͊;"{K��f�H�@u��2wA/�;��z�6	�d���혧`�{]c���I&?��J5ė�E��I>��.���r����΍ahq����Cy�E'̱�xGP̉����>i����!cG[��Uq!rB!0��*戹�*���Ҳʐ�V��رr�*Mj#�I���W1��:�iy�`Rl�UK�by��֐I��fMF�I�r���7�m�թ���Ԣ@�:Ss����:��%��?Q��jɣC6�,�b��)�b��<d6Q�WiA׶�W��[��"c���Rx�Ĺ�?�{R欗��-;�WU�,-���W����@{��t"f�V�7]��Ѿn����2依=��ږ�� w��pKz�VV�M n~�������>V�6[ħͼ*��/lYo�ԡ30�Ŏ-M[}Z�!�'rm���)z/�f�������TȀ ;t͏<����`7,
��e�ܹmܜ�1߭�����<�2x�|;���~U���V,�j�P�����3�$ˤX�c��!4ю�jev��*�����4.��� :u}��*���;.̂�6䦂��/ʞ�6H���>�|皟
$Ȧ/�bn�:ʜ��:��L��2��k�Ɛ`�~�'���O �*{���|+�����h~�Z~���A¸��!�^x�N�}�, pX3�?1�>ɀ|�t/`�vz��s����W���	d��@�"ޡ�]�UYH���[OHR��I��⡂8��THJ���!R �{�.PE����hs�%�t�K�X�y��!�VP�ؗ� U.q��Vu۩�=�
ZP��)~��%�kc5��ܸ�3\��X��G����s8�}�w���Pk&_�%�E�~I���NNN�T���Sa�FaV�)��>�Kj�@���:����H����8A�8��_%0�������˶ ���R���\��?��S����}2igU��	��?��K�uvX�/�y�'j�Ĩ�|��H�;K���+��҈�A�����&���VL��Q|��ҡ���]��o�b�,D:�j���`�T�?���W��rQ����d����mY�_�ì6�S���)���0�0SW��뫫_�ri��5�|�i};r�z*QIO�������v�+֬J���Pq�|U6pv����[�+Y
�0�����P�g"~�#�v�0Þ�fX4m5iO1�`^��[���n�Xd�)�x=#����L���_/��*@`��ǻa�Ϊ���ޞ�a^�:
�f�3��[$l����\�Ji^��,]���dMt��{�˫J��g`��%:�����:��8�@�gF]7"��c��xh�n"W��� ��}�G��^ù+˫��"�Y��p	�J��9�^ ��y������}��$o�
A�3�QYe��A𓸴NW��_u�d�`'_�s����� �
=��ӟ@\������9J�/�*�D�sdϴ�9�P1=?r1�k�rAA�D��׃E����ag(r�#����!�Xܥ�Оc�ը��_�iE�9�ҢJxF��:�vlQ_dp��l�C[�T,)$���F�,����[	GsH>�/�T�R2��%���a�79��A���.&�d\��ᩞ��=O�I��:qC�_!2�F��(�I2�qV�q��zZ������ TW)�e3-G<1+�V�d�ikֿ�n4:�fړ#�8���0Hp2��O����P��6��|.�}�ɜ�zs ��+�#+�#��rK�P(#�c5���%Q}G��F��Rs1���3�h�JZ��,;��̫W����Yє�M{�D�u��ϪE>��\�3]+�щP��+�'Nlt˟q䥅}a�Μ�a7T�]�GJUHuG�X ��Mz�Z�&Z��E��`��m�#���섩�I�K�*�Q􍓮K3��S��o��*�ܤ����I�Q�$X8��uG�y�w,���ϴPi���rR5[Y�Ꜭ���x�TwTd���A> �|ƪ���Ӯ�B�w���?b�d�;P��;Z��
˃�zy�*�X
��]�����`V	���,��皶�9.�a<nu^���}� �� 6Ѝj�qqq�;zy�vxAz"�e<�N#{���2
�H�����Ӱ��P	j�+�<CګM���T(`p	����n_ �a)��|"��VT�ƒ?�\��x��B����� ��Taʫ<dV�	q�f�/2�*�!V%�e��d}�Y/��� *��ɒJ��3�ˋ0#~й}��o5��]à_P�3Bx��1��j�]��=K+;�����X@"��!�J�	���k9��,t��`F�g���W��SIh��m �92�"���������Ǖ%��R��'+U	��m[`}H�*p[Ѣ�*�S�����T�JƄ�A�GT���G�"��^��}��M��]}�y`���@=�Ѕ#��G��"5�ei@�a�A���d�o�BbP�Y����,�	\C�HW�����'�AQgM"O�.�`N���(��\��D �+]~.�~w�_0ѯ|��d�`{��X
����aT�����Ɯ��
f��zG.�)5�oZgzW�3R�Yv����4-�#m����b@��\Ǖ|F�x
���v�=�l�?�H�NÈ>s;):$S��e�D��j�fO��\�D���@m��Y\GG�j6��JBL'AgMەW��emT��*�����t0 �i�����Ge�y/`֍�m��Pe+'�^Ǫa�{h�G��	!`[_6���%Z��@��N/�������-��kpGR��lU��`�n�lx�Z���/��W��*԰d;�μ��3(E"f�a������"Ff,>�E�a�o[�QصZ�.`���gF�	���qz����S��D>�#Яt�ݯ0=���U���j��o�M4Lg��@��☌�շ{5�=+*;�P�����9��o��K@i�Dl�rxNl����~uq~`��ZRM>Zc�L��9�ꅮ�0_�+��ܬ^�N������"��^C+��"��BEn�% �`�n���4X���YM\-!9]T�KF��?Q�D�j�.~#u��A# 䁴�\TrP�����RI�����`��2A.Dd�ΘCyN!*#,,�KKT6�3�w\���]�- gi��5"ՐW�Rk��o%j^!��6���������m�6�>�b�+���3Wj�l�@�۱�뭵?��^?� ,B��h���Q��tb~q3*��ٲ�
\�4&{��h���X)�H�t�JT�-u�h�$�����vt|~���ݹ�AWH91a�>n$��~�@\�����o��X�m"
��DſI+��}��;�aO��^x�`��U@?�I��ۧԚl��W���/7&h�Q��Lvzq�S�{�pZ�l�j9�]�)��zdSwQ��B(�	7R����":����W�*�	/��
��APS=�`)�P�Yl4]�cA�%�T��"���yZ���f���l�\j7�V��'�l��A���>���BZZ�A�0��K��w0SwC*P;��Lf;8��dMO�5DuzJXWx��~2��%1l ��~���=�b�(b��E�N���^�������PӏN�P�]�Θ]&�������#�k׮�r⮓π��c�$.~1���K�.�w�4p�#��O�f�l�Y��$�Q,��ɨ3�f��$�J?	��Ѩed��c8�]�k{{{���v=&�k�Ζ��?����>�p�T��J�/���;׃J��o{��� �Bd��լ�q�v1�Cd���Iim�J�6[�eY�<�Q<��-�b�N�}��s���аi����*&ƧP}����B2L�CI���ݺ�{��D�9! ��τD�����3E��	��fT�k�u����}WX���3RX6�'�H�~2�#������s�:���  KK����]��$.B�&�t`	��?l�8*PP�!D	=C1�S��t��D7���Vn�;)׽��"ĽeZ�<����>�����顐��^>��}��t�&� .mx���p���a�Lm�,iG6�F6j����;*����SJ�����' ���	��tU��o�b��˨'�/�m���k�>z���ն�U�]��Q���+!��f�C,ot<��{螘�G� ^� R;��@�n�yq
�
O�{�8}-��!����1C������fj��U�Ċ+q��-�����C�V�$`|�THxV���G_��h����V:�N)�ݲ��|��x>`�%��љ^�L�ӝ@/�<$ȍ5�҃`� QvȬ���5p�����y �9�VW�K\g��u��8]Xe��j^�o��S��@ǆ͟w�&�ο{����gZ�V34��Ds�6� z�;wrK����P_-��Rq>���p�b�२���R:��XQ�J���m�RQ������F����`Gb]B�����T>S{�Q��h��ÏpZ\0����R����L��O7��x��?}8�#�8�b�����N���C8�����D���c
��j܁���?u"���kѥ��.%<U:�/m$��y������o��?�M��<�ǠP���B��Tx2��蚘#���_d�RY�A=�� ��L���g�3L���}���T(_�t����~�5�����܈UJȈ�N��㶼rt���pSfXt�c��r5F�s��7~��~ ���j�4��Lf?V�##2���E���P�Ox渲ܴ��p��[���Rr?O�E@��S��Vߐ�sC[?BE|f��͖�a�^���_eA��Q��O5�o-]�z@�+IaB�X���.��n��Lo������(E��8��(ۍ��h�'��t�^LQ�e��'N��)q2b��C�ܟ�K���X�;+��디��M���>(�4�+��j�UtDP��6v$Q�l^���b�s�zo`���u��n�tJT�e �p����c��� �Fg���͍X@[�Ȇx�=<�y�l�3��.�^�b�9u2��K3���%��,���yc���ym�%NH|�(�+�ؙOB�,���x��:V6w��:��dc�LW��Hd�c���
Ԕ)�ho�G�IЭ���1�U��##�e�8�|������2lQ籨*�jX�ܦ�X�M��B�� <����{�N�9�Wو!�c�o����AF$�!~9��1�1!���vz3.e�4o���N�6���EPU�3x#�#�����cJ�	�rD�����S��E�$_���d�>���߉�3��k7�(��uэ��D��b�9�4?�*�:���d���! U���'��b̏����`���
�%d,--O�I9�5^�F���v�ޓH( ���o�>T�n�����TYZ����h;�32o�����aM�j���{�S���,�&��3{�p�%��� �l�����O͙�m�j���=�c�t����5�a=�,�Ļ27s$)@߉(����E��ag0.�@�������بc糬;ZX���mo�W%li�D.��s��[�C�Cݱ/�$�;ܳm�l�U����q`J����W��������UR�HC�Q����/�e+�}q<� �W��m�Q~N�U��X����P�9"*;^�Z�c���#��OU��6�ӨC*ܶ�N���¼l�f�2����6�; P��A�PC��`77�����%�@�L�IÖ��@ �z�ԡ�.�xk�M�c�Jm�K}X����CҀ�a�>���7~	��b%�q[��&�m����bv�F��;��vgq�&u�<��+�0�L�J� 9��e��i��o�C䨙�an�I��ڹX�.��:���E��N��,��6:A��'�k	96�9b�:>�ժ��g�8M;wX]B݄8����*gM����3��t|8_axLuR1��JbC~H<�Î[��S�&�=������7�I.��~E�M�O�Kҩ��qQ��C�m�Qi��_���]ѡ�i���#�`l���|�.����V�P"�3�̛�z��^7d� ���$ v�f�m�~�\W�~�e�3��]!�հ�]K#@U�U�>g��N͏�� �o��v�p$"m .��q#�76G���A�g6(_�l_�4�.X�֕��Nv]�JBuC���?�N0�^}+���V��9�ٗ��g�u1��oXO0A��W�s�?U0���(B�u(*%5U���&ԡOܢ����f���:�Z�A��u�C�(2��K��x+,�5�&�>�Z;�|L�X?0��_���U�v!F�X�\H���8.�qj��-�B�B9.�HZ��.tq��S�ڂv�k_���'�?;G[vĬ8d=��ܹ
c ���$w/��O�zN�>�l���y�LP��+BJV��ٶ���Hݎ���d洚��#��6�x��6�m���^����3��!v2��P��EW;�D侳�x[�x���9��)�j/=��h����'4�a4qy�-|��nk��ßSCO�3��1�8#q(Q���{��0�`��D�B�Q�^R�b'u�|md"�*�n��6���A1M@�O |�#AC�Ųݞ䫇�4U��{�_�ӧO��Z4h�Ȩ�ԉ���џ�I�t�ۇ'Z�uʉԞ!�b@���Η�������h$���O+%F�j��M��F�'q�D�F��򀗄��;Z��~���ܬ�: h��w��Ϳ#i:��F��5�F�+�u�j�,��ǌ�q�^<��	Gp��b����:Z�>j��C�S$#���q��>~�Y{���~����-�=��;w`y7څdo^{u����`fF�o��tbJ�Ψs�V?��R��R�Fi����yԞ�A!�)��%���E෡��"k����iw $���
�pd ����w{*	��+�<<w��^Β�Ld2�_�L��e���y�L�v�/�Y]��	˖�R ���hy+�m�J*�3ˎ�N��o��5콳�E��m\��:����K�7
�>V�6("�d� �J_�U)o^�f}��ia�.'�~��(�;w��91Y��ڧ팑c��6��T�-,���~ZV�|�h�9�F��S���D��*u7L�~���o�NI-�iP~I��B���G`�Xs�2���_w�x[CK���X*
?"A�#L��r��%S+�.@���@����+��M�<@aޠ���"�w�(v3�Өٙ�)��}�[.��$޳�3�
�tՀ��s%҉\�QK��T�4���U��d��TJE������X����Xq���:OA�q�A>#��a}'�����n�rN돎�5�7�S�t��K�`�����9yO�ׄsވ�`�)ٴt�q�lQ׮:��b��O4�m
9�������l�U�Aw�р*��t �����N���7`�Z����,�
NyO��u<���`f�۵��~��'d#�ws�w;<'�P�
��8�o����-�d�8��K������޽��������� .�/�ϘtTΆ1�Z���5Ң�,e����젎h ��>������(�p����F���zh��~t�i �"����������p�xU�����ml>DA`2�D0A��C��m�;���0ӯ��^كZ��W%��R����Z��OqOzZ�׿V�|�J\���Z���<�m�#�vK�?�N:8揎0kD�^�A*��!�%Q�?LN���{�1pN��.&� ��Y��j��,[L���B|��+S��Αu�d~y��1r,���z -	xdc��4L���H8�]�Ī(�&���k�m&�E�!K1���ذv�O���|?R�a\�x�l}jξ�;K�Xw�[�{�3툧�D�.?L5���������}���"����c*~j��r|C��E)9v����M�
����q��MmQ���[����!����ne-�������-��SAqea��站��<��ۙы�����P���4d\���_�ol<�y1Z�������b"�%]=�
وnƿ�K����x�Nf�u�~$�,3:���e�9�X:҄�{�J)��yC�z8�ͺ�K�XO�[=�^�������/2�;�:�D�1g��!Y��a�8<�j˿ՔM��Kxy��1m֋Ԋ����-���N%�'��S/�)������@�w�nǹA����sU��6L��6��~ԃ��m�/x��ۣ���@m�N��S���/U�����la,�'F1~5���nA�X����.Q�������{� �KA�U�sd��;�܅��@���xDM�q$�7o�*1��yᾛ�O��`bo��d�`s�I�ܥi�o���[��k{��]F7��,�g+&��?R�+���� ������� �A�X�a�7)&Ǯ,N���a5k�$<�6wu�q�3�3�����Vvz-�z��;�t�>���n�c�0ٴ��c'ԛ?�a�,��(�����G�tT�z�AB�ɸ���%L�'��R���%S���C�%�ǜ1�i�(���������6�����c��p����]@=>�Ÿ冲cE�T�Ie�7t�?(��0LEy���[#j��zN+k�K���[q'�MC(����?��������]�Y��Qx���S�j����<��p�梕9�f�� B� ���K���4.C� ؾ�	�2��{c&T^�{�kyaR(��'$]GW�)�)%Ȋ�C�d�`bY���c�$��}`�R,-��������Zv!?��^D/� ��-�r�ڣ���-��"���q���X|%j�.!H͂lzt��/je�o��400�����:$'GdU]ǯ�B��XS�:Z������"t�h�=��aqv��2�*x���3�Ti%�[��]
�z��UWn^^mfS�-֧��G;,WTT4m��;���S��sP����}D���
|���K�{_�s����X����2m��D��5�]B�)IѦU+c���l�B�U���	-%�G{J��}_�uݟ���u�;��:���<��x>�z��u�o�(v;쫌NH�s����A%0�x���)����t>Rń%0�B����	��������o�uvLo�����v@�����!b�]-�,9�6;����`��d�Js�n��k�u5%�e�3}W=fg��Jص�w*u���N�9�9�軿�x�@��� �k�,絳i�%VV�Y���=Qe#��0ծ�X���J�^�BG�|��ϯ�0�(ɛ]��>=1f�/0�d�V�G�gǕ�N��6Ɓ<V�}���p�,^�f��YM���Xcw�ga�Ի�=::t1Ci�j�y�cRX>:5զ�G����<�Hu���T	'D��8W�|sr$�Ư��bS$y"�P2���V,����f4<fG=�H
��-��m���T(ۄ݂#�����
K:ĚG<=g�'�V��a�6���� �F�s_x�['�wI�}m�8?�2^�+>`
��]�5t0嚖��sp ��_����%�q���j��N}�]O����0@o�h*,�9m^+�aA^��Gs'�� o߀�c�ܛ/\?Fȇ��o>YvZH������?��D��Z�����+ ��ڴ��BERI4�xP�)+�tù�9/���U�K����&�6ݭ3��d`݀E-?�@H�k�"������ةkiF�b�+��"�Q'�랞�=����d�[�(�[��U\�kT�ho?�}��}6�x�Q���?L��@���%aͿIMj}���p�����43.L��C�����>�h�-���RL'�i�����T�MӼ{�z]³E��5�v��2*
��@�)@̒��[X���֏�'y�F8�T��<8��=�)����hp�I��7
��]{n7�N�2�䊠#�`�bՇ|�,�5�k��lf�\���9�ۖ�sc=?��$-e4�H��e{����e6_
vj).��Df;�r:66�fo�lo��QtwEo�>���Gp	ƚ�i<���	�nEc[� ��a���S����7ÒKTE��xv�eَ�Z��
-�w�y���(���Lo�PZ�5�`����ɒ��%�-�#������-���c����J�d�'G������T`T��>o�u��I�Y�/?)cb��B;�VN�n���^��%=.�=�TC�����u�Bc
�w�D�.�������t	*A��PR��(=�;;M3�M��
����iV<x�߻���Y���	+�{,��2�϶���;l��k�.T�*��C/�tf2����8��[��GY�X��<rN�[�V �t�6�d4$xs�.�ݱs�\�85��м��DlĜ-X��ku��Ңb,}р����+�1���/O�����X^�M˗��}������~%U"�����8��!����[b��b�7w�ĐP�h�ƸNw����,sk���ak��s�-w����du1hg	0�$��)&En��W���Y�����]K�VaP��2�YЋ#�UL��<��l�p�O1��[���^�?Tpa�iRqHE���4+{���߇�]ad��]��O�����(0Eg��� �ws��?��H6��Ec�K���J�����p��.����.]��bq��e���w��X���{��b�
��S@Z�.r�o�n��m 8y�/ɍ?C�/ ����l*Bh��u�5�Sv����?/:GE$a���� ���JhT#,��]IQ�;�G���������-'U�`���c��PCׅ���d�'��/AF�
Y�F��\�q�3��v^�ӏ (g�
����^�zjR|{�Ý;=E��:=-~=�6�[6r�X�
�aAᩞ�t�;`K �G��g��*
�������n���ŏ��3��!-H�y.ͭ�\[:&���1�6����w�ӹٜɞbF���[�E��|��>1��g��5�L��Z�0��Gj&�4�P�N@�_Ϳ��?�s	�5�!����|�Zʳ��	G���O��Fv  f���R�^JII�u�V|�,�>,��������ʭ�u�A��LW����A��h)���?�}���ݗ;�N�����"\EY�����2�O��4Â�jT��$̑%_H���Ę+FK�o,����wqq�h�.�5GU��~�|�m��S��/�w���n苙L��~�?�ﵢ_�cX����j�`�#�S!�yE�#��1�>Ăn�h��U�ww����u��π[�r*�"�շ�a�]&�"�����Y������e�������o�
 =����Xה5XR\�h/��
'���: �R~�q����A3�D�L=וX�T
���_u6�N/�r�zޗ�q`� �yay%��)4��yHfN��+��"��n�$�jTѥ��M���4d����D�����2����n�l�6�>]��s� %
W�)-��w&����;g��ՍE�a�H��BP_/_�� )k� �n����������/SB`|�ܩF�R�1bDy�ݿ�鮫�o@�>˴�J�HW7�t�R��g���)���pv���^&IQ�J����̛�0���++W�֞=���T��YEĨ�8�P��٬s&Y�x%;� <��/\�1fk2�h>�ȹ�;S��*�>�:��~n�~nD���c�����*b�5�U�V\G���b�j��|�y�`fn^����J�y��aO��]��D�'�ݦ���(u���)0�
�F{��bf���\���D����R���K [�b��K��h�#��k�5Co��s����������؂�v�-^9̉����	����8���d/&��i��D	��Zc�;:hTvq)�`B���ue�����65�N�-�j���OƉ5)]޻��?���ij�'X4��'��F��a�����;C��w/�Rb���/G���>�ҳ����_1s^y=��9�ȁ�+��d�C8���qFs���h%����_Q����������4�6�<� E�@��K�ZOVc�̏R1����NRY�b^l8�H2f�Q� �fB�v�E0�]����F���G�	41Μ�*��~ z���{$i�y��Ɲ1E0�g�D�x�u
.+�IY@�rd��ځ�����gX��"��%+�Н9�ҍ��rr\i����(��kZ���p2z{��h�=X�$ɀ��[\��D�B�<<F4Y�b��r�P	��1v�6v�kLJ
����_䤝�M%�=P���cYN6��[3맅 SoB�-��8$d��6�����UQ�o��+i�GH�2 
���%2��e5i6�S�����[O�z�IQ��-��������F������Æ���y>$�Yc=��c�;��;d�tH��C��],OvI���~+�.o�`h
uE���4�'á,4���X����S�爋�ѷ�� /�F 0G���3�u��^|y㏠V�Y�Oi��4c�H)k�9^�;��|�͊�`f�- H6�RH��W� ��E�\��M��`|n��K��ɺ�?�I�5��O;�Dq�g��_[+{�P�54�l�}��ŵ5����mѶ�q		~$�*@�wV�!��j�!+�~��Ѱ�|v�6C'܆�����p�2CG��J�4Ao�ƽ-&�kƸ���u�?�)��w� �V�8�;s�n�#����@��M���ٕ�u@����#��i;w�,�&�ob�f�����$!��M�(V���֨)�j�ȥ{r��b�b�vh����ѫ��v�5�*��c�c  TA��L��Uű����"gZ��1^�/����ƣI���%C��<ͮ�ʏ����E���S5����B򅞙z��͇_�!w`��b�#�4y����B��AAAԨ'����9�f^:��@���h���_qS�Z�[�1N�1�AB�Qh���)=��
��W�}�Ġ������F������2胎ֻX!j 	�>�D��ִvW�e;���s�Fr���#p=Iʹ��X���߹w�0��ޗǩ���w���t����L͑UG\̦�����Ȫu�#@ʘ���`�:�
/�jnf&R�����ո�{����v�f9IP�Bө:�4s��]��z8��
,WA �[.|����diV���"�xkt�s�u� ���i�k8���ze�:	]/�(�K]Ĺ!��p�zna�Y<�ӌ�1A ��B���/�o311ѕ��
��ɿ�]8=� �w��c2HH�4�� ��}�A��Z�%,���:s�(�Ȋǭ����f��	�ˬ�]6x�h�����P@�J�h�g�1 �����.��$�HU���߯�����,8�����\V;9�͇�j@Q�0���BT��w���D�.Rq�lj(R��4��������p��{ ����k�����D�
:�96����#���&J2�4ﶶ��7*`��i>9�(�s�)`�&q&�r��+z5n�Z�n���o.�������=�kb��ps�&q8�W�8�����x�(�Bȭ��]�����U"R���;@�|G�ʇm���T���Xh8����U�!�X"�a�'%q�7��G�{�������s3-�C�Nz�����VJ'�����~�,emG���@*!A�ZE۬=F�LXqN:�Y��c!2HOD��c�&k��	������*��e����.>���	M,�G���+�fU��C��M]�j�N�>e��_�͉��0o��n�0ֈ2�ѥ��v�D�w^��؁�`��ڴl��z�SÔ1��.�4SS���ڬ��>�X�GK��@�ڵ��#>2����@�t�X��) > �m^]�����$�L�q� ;^?Sϸ��&�hk��bx���8�v�\�����	=��$ʋ�>�d8����$�R�FRJ.	|�a�:�ũ��:ߓb5��<�o�ϐ��@9���@�T�C�)��v�I�?r��7�9�{�m�sㅅ$��{��z�"�&Y�\E����_����G�N��Z��L�߹�tUq�#Mjj^�2�C�Ejr؜��.��zk��:�eO�MC4(���͟i
@̄bRq�&�.���&X�F���ن�q�xX4��g�#��bf�t���.֑7Z�)�쓔iɃ��Q%���saL� )b�^SPdl��4��U���
Lҏ��;�gW���W;k��]��C��f-5�R�Mox�ڪ*^�lsް��";b���ܢ�B�n�������*^�o@p����k�LP��^%%%R��>j�v`��&hR�CM�qE˹pP��4����2�ۚdj��E~*EjZ&14��Yg3������%oT�kIi-[�y��
�|������ϋ(���))$��E�ԧ��c_t	C?f��9���$Ji�&E/)Q
㻓�O���Xl�{a�ʹ +"I?V@������&�N4�|�O�.�A��@ ���IrR����D�^꤂A*� ���(^��T~X�|#D��:��L��rD�U%�`[)�$�0g�諽<R�a��`��M�������mF=���r;Ek*;�:ͦ9IBԀ$2=$���Ø��ν'�P�X�<}�zIp	��$��0��S7qyψ
�~�
��D� ���}XՈ�G���Z��{a�'��fVV~��НY�����(��e|M�nx�.t;��)X���@6�v���9K�Hp�J�{����J�U�:Ds���(/��̣�	w�o�־3�QThYm����GMR��#���Qdm��;	$�s���_(X�z�X3��dz[0B��Dm7���Q��H��}^��,P��od��"F�{�5C��@$C�(ap�}I� W�vJ�U��&�} �ۜe+c�7��P �H���Z��h\�1s�N��5�f����朱&r��/��*��Q]��JL��/~�>A��̇1 ����@w=;���$����a��:H�gz�P��߇Z���,�*�$+�ڈմ���)6,������D��O��'*v���A��N0�w��׺_� �K�`5�*-ޯ��o��l$כ�.���=��
U".}���}ٲeT�a8TUM}e����̮$�h�`D������;�UЉ��Ō>eZF-tl��G��OG5ͽ����.0>�z�J�#4��T��������1.6�K�Q'���a#O��ы�����tĳJLL����ğ/�K�sz� � ��}��M�v�����vf]��*yg�����1}�t��Km�<�(��A\��F��,-�H2���>}:�]�"���L{�ɾ�?���忘Qn�Ҹ��NH�Y���,�U��t�-����*5�E8��vw�:�?$�`�-+�DQ�B�⊁�!I�\��$�>�n�tޢīV�AT.$}�����??�|y}�`Ѩ NC���)�I%{��m�	�U{{8l K���o� .���b�G|�/vZPU�+&}�		��?��m%]K�9L�~R�b��� ���R�X�O����dT'�}��bi�+7������$��X�^H�Xk�,��H��R�V���M����������L�ъ�0,���^��U`J5����FL��R��Q�a=��N?���N�oO!0��� ����-@pr&}6Q�#vӣ�x`$uv�)k0���� Zؖd��d�H�<���ݔ@��Lğp-J/��B~;aR�q����+���I�oٜl��g�ja����ߔ���Gн�>qi�M}6$�?�;�Zj��1��\Q��k�9 �/I9s��&U�+�coM�fh��^d��Dl�����f��ڍi�g�4�E�4w��F0�����Ԍ_��T���L��8C�M2.˃FB�}�}����gb�ňTa1x����������5w�EH��R����\⴩��~'�Ay��Wz�&�d?Au�����ƴ�xP�x��:��iJ���������X��JJT6�F�fn%��/���؈�t�4�~|,\����ǊL���Γ�P��?��c�Y��5���;bb��s/����?]x9��_�:ijw�X�_�5_�d���>w+x��Hf�5B.!@�ҿ0[�d�
�ӓW�,�+�<�]�p�%(��;�f=)��~ɫ��`��/�Sy�ޯ �aA8�7IM�n	a��0�k�^]a�T�J��#��D@�	n�ձ8�G늆��NR�.#���,q�r\ϭ�s�";O���� ��k&��N�����a�+��,�d��e�Iu�qS�?���ڀ��Ɇ���g���%� �T�`�!�T.�:�n� l�4�-��е�
��OO�t�)�<��ĊV�Bq���F��f݉YDL��痗0s�ki�Ϡ��y9�8�`�6��no��|r����c'ô�n��u�q��2�eZ�H]��k���N���8��Zj�H��Aatd�*��;@���5�V����I^^+���R�{�	�Q�bt���Q	�V��� V����V������ټ������k+���������b�6������a���AT��LUTBBB�c�pq�4���%�J�T?<ʸ�B�+
A���k����$ \��o���:���0Y�?�1[Lv]��cݭ �q���A� �aʝ��0�@RaR��1IA�"��NX߇�0X3;��I׿�0f�5	�ϓ��%�	~���c��T�NY�c/�C���W��N�Ǯ@SW�����)O�h��hc�j)�=��Eʽ����z���6�Kk�T�|||�x�-K��+1</@.!�h:	�JCJU�"��E�f�� �8��m���40Q��7!���1��S�ͯo�cҔ<y���]M��U��Yk[*O.�~����m�M�Ci�&9��$b��xGK�2�B$%%�B�� �r:�(�� �3z_�eJ��yI�|�M�C���������m��L�Qe�6�Y%�i�&p�@�N�LP��V��)�)g��"J(��666�p����^	��YY�nkJ���
}x��%�n��C_�[3�jk�a������134}�?w�	ӝ�Į�n`����`�ПEC�<��gB������x:I�F�)%��Y8_Q�@:i�tŰ�����|.3��9�8��̙��A��NI���C�-�gε����4��r>��y������l,��w41}�7X�4�܄Gp�k����]�[�"�W`tj���!([A�
�(�������!DXwjCp��J;bF
�`�l��8�9����%��XW���^@���\0�!��߮�o�œZ��:����с�o�oT�w���a�A��ra��𾎩ƑA�
�D���9��3mjS�=��ȿ��%�⽚>>~?KP��31�mn�����Q N���4����t�Lue�﫱	92��*1c��/�k-'�}~��_1ƴt��-x���ԛO�?D��&8�O���}�<���wfH]�6x6�I���Ys�y���?�9�e�w��9�Al��
�~�2}ss=}'�%�U8?7{)�A��)�PM�I�,3|e{^�R��*�=�!�vG� d`��^�cv�J��G��5@������88��rAGڗck�z��;%77�ٲV�,^�`t�gA[��;�Fp�`�A7b����&�;U�8��Q%��+�y^"�T|�@ Չ��7/�Boo�I|��G|f�F�i)/>�Z/��FyѢ//�V�Jje��'����\����s�7��n�1�4�h�x�}xo�m�GS��N5���s�(�߼?kWj���_Υ��K��V���������{0;tމ-d�VMM�D����2a_o֦FDl��VR~��a�
��'JH���	_p�����X>�TZ s�.��j�����/@���.~��̋�7(ʌ!�0;�]0��Q�J%�F-�	l�r��O'��GGDDD�����׬�i^F��Y��kD�6���c�J��M�U����-�� �[-�l���~�%�s�a�wL^�C_�u�l=�R�ǡ'U�L��\-%%�uS��]^���گDj��o��/���vy��x�̦����ێ 򳅮�d�LO���?����?�f�Ut����"`A7�ď&��	P�FW�U�PA��FԦDGG_ś@D4���&8-��"3/������Ǥ�~C������VWWk28�w�Ύ�)N�!l���]
!~ڱ��aW��F��	�ˀ�&c4;D�D���r���: ���%�����fj���W=�]�f>���NJ&D�AQ����R��F	��nJ|�:wơ����������1Sz�\|i����Ҥ���ZX��ط������kl���7�䝊4�f��x���m�Dh���t��p4>��tl`һ�­�`���*��g��	����oa[�;b
Fi���;�؁�����}7H�f���=747�9�0ݮ/�x6ô����1�Th��76�X�8�Gs��W�7�F�Op�wE|�o�x'SL�
�Q�Gk����S͂�%l����L׏�H���+;L�XfƝ�����v��3�}��捕?b����w�����=uJ�~A��@���_9H��&��J<A�27�J~���ÞaA����`~�4y�3/`N�`��X5��s�wK�hs�H'���{�K��-[���Q��x��R;t�X95��;
�U2>�֌�H�
#�ќ�1��������ӛO:�wjm<�W�/}���}�zL�jE���@���mX�/õ�]� ��k0����O�'���~�8�!�_s�Q���,��<¢��A7��Iw�����Ԫ[r'�-�ކ(���*��}�� ���Z�:A���+�u��d��J$ɽ
!j�C��f�j���� 4��E�{��{���-�L�I/��DV�)ǒ�YS��z]��̭�����ӯ���ZB_"#�n�AaV�>�}H;��ЧJT�����1�a{>���������7���|Wt;�%�7���2���&ø��%f���Xd��7�`nU�3/�m��`Gg>=��Z8G~{�����8��5&�FQ+!��;�ϙ"��� ���#�bW���r2��Z��}Eh]��paz�#e�7"D�2�/HaR�C��D����xx<i��iџ�B~�HK?2o���/鉝Ɨ\���L�An<A10��0;^�*�DM�����c��z��_�zj���??a��X�j�偣>h&�f��t(����;�
��������c��=���K���?�`Dn���J�z3oTY�sM�qU��7c�����#���x�{<��������~/E��<�y�a��2�ߌ!���덄�ob�>�<��Q�^��<C2��Uy�&'Km6Ⱥ+�{���0������L���;�v=��<�g��������X��i�) ����,�ۆ�}���Bǰ�w=�Q�֫��L�?�1���$#}�\l�����������%�F���-Rъ�JFK�_[�hjy�nJ?mFY�|i^��g��1y+�m>Ǝoզ��LbQ'tT���9�p�|�ҥ�U�zv(HW�L��ȧjA2R'K������C�ŗ���=E�s?�!�L��ʑ,�ڳ:$a� zh2�/��̴����񫊊Jo�=p>�=���Te��s�pz�un=�~<P���&f ���>VF!$�0��Rt=۪|d��Y�vu��N|^����!�d�ôq��K�k������0r�r�U�����ʹ(z(��+����cl�lB��=�C�VHS��l\��n�Up
N�+�
;�V�L���o�	5����"�p��X�4���$�	�tU������8�7��/�����t^�G$����~9�N�'e��o��-5��WTTDm��p��"K"���+�m�8�8.�7�\�U�*B�41a�`�?��1o�<|�Bd���O��U�8l���
a���TЭ�yn���+���g��k_�R���*
���[w��zKuM%��w�pRY��p����ş���3{��b���Q�ZB��X�w�]�g���p.����
ȫ�OS��k)u�o���cN�ܒ������������W"`���= 2$EhBj��~�} �����CRR�H�
��Yqm��`~Z�W�Wo��	C���w_�	�LLZ���`���1����mƃ���'i���Z^�k^b�ׯ��6���OL��?2yȄD��KKz�LA�
�P�7<<m+z~�/cw���p�^|iJ{0n53zeS��UR$1[�7�Y�p�]=�cP�����h$)Ju�L�}�7����L�p�ߴ�=��V9��_۷��ֶ���&���NL���,!i���D��Lw6GG+�p�5H|�8���qG�6�rN��	jf��Joo0�O�>}�Qp ��ŇA�q�z�"P��a|�)�w�������z�H�0�b �7-gWH[� I���]64̰��3��z,g������K!V?�� l|�~�ky��P���٨i�t=a�;�U+���o��n�pd~z�!ز�>|ϵ#����3��&�L���Ejd�zR��TYY��9©u�X�ZVV�`�n{o�ZP�8�鱎�j��*�OE� �l,��p'��D���5@�}��+f6kFrU�띊3͊�-� \�.N�[%����5S�%���QaM#5V~��H��!B)�8�&��C���=Ht~́�WQ�V�፫���mx%�/A/X�@3���^[�g3o����@��PaY�������in�I�	�
j�cυ1��E�]�a�6???I3�Y��'))��5Vo�k&��F?s���"��/?�j2�SWV^�)q��_A���LK}/_�l8nk��U/e�oƨ�.I�|��v
}����UO��=z3�-8 (//U��E�d]�o�m[h��ۺ�W����E�����1!��6�9���.��E*Ʉ���|�i��O���5fziֿ�+
�z�h�u'�>%"�� ��B`4��+�������7�B��#��>�ٷA��B��=~3�|�զ�m4_,!�&��t��Gz8f]�M��׊u�5q���I�?�G�~ML�/f�\�~aYe劺�:�6nw�:��Dp�W�N�(m�\�]�����ש�О�ύ(l�ٝ�ĕ����X��s#�FF"T(z�������U!�� V��oEEH~�R�k�W�Z����N�M�S��f0�l@�wv^���i���ъT՟}����'<�V��Y���a����A��qw�w��L���i�'�|i/����D��(ni���vM�q�`t��%a4T��-_���9�%�K@��V��ǿ�BJ� ��ޓ���z3��@��ں�>#u��{����#�˛]^�|{w��DȞ��}��$>�$��FS�_��*Jݪߕ;7.=��a�acQ�!��e��N��V��J�d���_����E�~{�P6�HĪ�
]�EL�����}�B��$aQ����d�����\�(��}��gO8�`�pҹJssw"�,S�TQ!�׳�s�A�"��>ԇ�ǎ[{���I�+��5�-�K�Q���`g�`ׁ7p*�d�*�sڂPD2�љ���"�3������[�� ����*���ӕe�?��bs�ͧ��6���7�h\�������=���_Ǚ
v��Y�eL0��zV
��鞘U-�ĩ���v ݧ-Ÿ���3�k�㏽9����jD��<���@c��{�_:��Gl䩛��Ӝ���$��0NN�+��!�B���eT�'臏�c_2�O�Q4����Rs�_a�c�E���l�O~,��Ϝ��w⌋�#5�����Ok֮�{'���f��짮U�ߴ���r��l8���Y_�|�,���i>uqA��#�,��X!�f�:J��WPQ@<g��ʨ��Y���~!�!L��ǀ�B[��P6x={���T�6����(;g��6�Ź	�ш)P�Pc��?D}��j	�%#0bg|�wͅ$#���p�(㙄����P�aأ;��,�|�'�<פ*�ƘP��؝��M�qףd@]�/��[��2?5������I	/�:���A"A�H ���`a~
�\���.F�L�<��ŅL���Z�փ$i�&cpmP�U�`ۋ����q{e�*p��6�������ͽ���}[�SӢf��Gd7��T�2"�s��bY��)�w*�������ǻw���qI"����^o�)FP�ŋN_#��V[�!do��$�.���Y�1\����I�����an�����Ltx�|���!߂9ɕ�X��Sya�B0-��`���=�����G�y��%�.&rc�� 5�����SV�"=ommeNK��@j�����h-���֟w!e��Z!�"V]�Bd�m�vV�wuyc>n��a�K~x�ٴ�`� ,��[Lv�D=^�wW'��Y��	�*�ӹA��i� �ga!ݰb�%t���iҴ���foX���>4�"K�_I����c����>��a�t�����hT	�>��_)*��o}}=���@j�-��A���
~�)�����r�T�,e��ѽ��E�'6�!�~o�k�yl�`łL,Ȳsp�(�!�����/������xˇO��#+�Y�h�b���`*z�u����$2�ϔc@��0�˰Ot�Ǐ⨣D�{��F����0�@%uw�~���EI��h������u��={��̿'a:'H�Ѽ0̋[� M ��T94_�8�X?u���pU���o$:���3�X��������ZB?��,�?^�!��U�W{�#�<E)�һ6��AR��������b�4C���z�j�����}q8��`���à4�0��9-�ĵ��x,��H
�nC7�%��Z�<���L�ʆ�.ED��	�Z�ti޳R��LUgN�Ɲ�;���D�:uꯠ]Y#է1��.��1H%?6.������_-�����F�+��ԘFVYE���J٧O���rPA�-���x(0�P`����1��ѱ�P<SL�����
ڶ�� 
����`����Qc�8&������B�ۀ6	j�H���Y�;L�`6�2�;�G�ӱl��L�cӈO��g�����rr���@��J������ѩ�Q2ߛEm���)ժ!�5����@$w�L@\!�q�o����]��򮇿$�L�c-���0��;����wj���Ԭ�d����*!:������Bh�c�����R��̦;��o��ݰ���;���k���RS��?�*U��x�Ԃ��Ʈr
�)�,��1&�����28�ڷ��'�� ��7�R�0|�]�r�����&?�(�t�6{5>�f8:���^*���K[I�5 'O8�|��u�믉�%y���24]�<�(��3�u� ����� ���k1��ly*s�/���G꺈��q��s�����q֧�OY��>e}��������)vU'�_r�xt�u	����;˃�b�X�����mb��w���j�Z���j�Z���j�Z���j�Ok�}���q]5c%*9b�?߇�X-V��b�X-V��b�X-V��b�X-V��b����2�����o3/V��b�~�t؈���y��׺o�x��X-V��b�X-V��b�X-V��b�X-V��b�X-V�rk�C7yL��uڰ���5���8Y-V��b�X-V��b�X-V��
����w� �m��j�Z���j�Z����J<]HЉ/N�E&�m����+�;~�)��j�Z���j�Z���j�Z���j�Z���j��lї������~_½5��Ĺ�������c.Z��׿.����;��)jm������������������b��5�����>~��?|��Y�d��5 k@ր�Y�d��5����kzz���م��5��*�ږ�Kt|��k��<�f?��+ެ���!��.N��]k����94���[}�缸(�ߒ�����������Xqa卤���lO�iK�y�+)Ŕ�Y�+gP�}z���g�{���I:�mZ02�E����u�.��f%ۧ�E�GJ��&KO�5~�a��I����O��Jac�0�۞�O�^F򎰓Om�έ�GW��|v~.s��ۤ0���r��&!8��z��:���-EI����coO��9���c�.r�8E�����e�ů?Q-��x9�����E�F�=��>s��&^"�����cs�������:�\�����l��u���x�H[k��F�f�V/N؋VT�z����1��_���X�7��0/�͉3=חYԴ�2���D��X�����j�������lΪ<X��8r����6_��r戡ai��O��ZTӂ�lmm_�)��w��,�z��tS�y.����̝��q�ec�=OՌ�o��>?�����N|�t�����%��$�a:�t��ٸy��~����>7�_���HW7�k�� M�;ǂg;>�R�Т��7�ו��46����̭8y�^�/�%i�Iod�@~�-�W��E�5nc�M��$o�Rt+�u�l��i�A����jV��:g�K|9V$�m��� R?~l�L�.��/��;�� �o���F�;g6��-�ӧ�'>~�������
�m��)�[��L�2�~�&==]&\�A���'=!>�U���Gt���yڸ�٣�����׀p���Όq��J#:3�;���ڿ}!,�f�y�\'�VK?����t>�a��3�ڕ��W�mH�5��[J��Ţ���O~�ٕ�
[��G�pv
�	�͖z�t���$�ky������b��}ʀ�{��v�G:�6���_��^�{�d��B��7)�m^����f?E����k)�ms<�olf&R�(��I7۫�*��x]m|H����N�뺉6����]/^��Ñ��Φ���،tU�Kv������K�����2��.J�x������	�T�Ġf_�G�^�G�3�}ԙq�������\ⴹE��k��+3kA�]/�P�V��Z����@��>����^J�nW�|���xk�ۄ�YSa7�>}S+9+�E=7#�]��	U?�[��;�u�6��{�+2��c^����;�-řF��11��H��;��J��QHk^���3#ͩ�Hn�=̦�6���nq�|F��p
͵�6C_��9֥ɇW�t��ON���4�O�q��N����}��6����@S�j:v�����+��efw�E�B�#l-�Ͼt	F�i?M�����fI8�kz������4ڞ����NjKuixCo!t�����ʫ�Gw9$�e�?��Q���o�Ro�dKB&��o�O�N�iJ���q��)zy�O�>m�y��ѫ�=,��,}��k���V���A�Ӎ��w�5���� ���କ��=fݍ��sMlF|s�-1��T�6ǒ��.�9��!��_Djɒ%�[����t�4Z�^�8��у**ð��IfJ��;zG'���
>b�O�n}zbRүbbbt{��c�k��-GYK4,����N�h������`[�Ao�#a#777zNK�e�ԇ�6_?��;'Z5�|J�2�1�jp�2F8���Mv8�^ͻZ�k/Gyy���	w���������Gdm,��T|#1���mw��}��;&��{�;̓��T@֯2�%''��p�wg_,
1��IIK{�x#�������Z%SSS��Zm�jj�������V���ݹȴZZZ0�����t̳_$��d��d�}a���Z���=���L+�k��G���?�`r4G�� ��ɑ�k��çj�)���4!�6g����F��2������8{5�󄄄��`���c���읾5�ւ/\�~hܓ����C��D|S���O��*�}��mm>4�T�L�>yy~��V�ϴ���oLA}KS��IB��o��j��WY�h��t��u@'��`�l�!ضQAQqv,ѸP���pL,M4&ԧ_����w�;�LL�>|xmӁ���4��/���6iUf�ո/ق/�L�U��_�:�[Z�,��u��o٧j����S
���1j�qۺ��Y�&��e�5�i� �<i�q���w��i�O��b��;�C�u��I��*�>*y>]k2�u�BBf��_}nx�lYm[[��sק�%��n��O���+�׺�u�#�`�wZ��y$����kv�f��#_36wd���I�ګOO�A��m�l���	ǵ/5��'w�^ �P�J_ۤO���)����͈�^AW�K�b&G?.&�g����C��S���x�Og��K��<���C�}��˫���W�g�ߢ��i��>�笞>}6I�k��t���>�L�������'���t�G�11��\h5>Y���m:��^%�c�jI{��:�[%&�2���c��;�7P�w���i�3�:~��#bbr���{
bm'�sN��q�
l-��ˑ8�86�Sth	�s]�p.�������e��b^F��}�˛��5�<	��Z%[�P�����G�6��}���c��=��r�Z�M�Kݥ@Z����-��
F<I�*�5�'�j���0[	�I��I��0���t+L��=��w���q{�/<�Y�jn��I������P�\��g��ٔ�ՠ�穕kV��r�2{����I�^�,�֞n��F�[��3�E�t5�Z�ͼ���N��/>�{t
�J�)����Ŷ��������I��2��O�4����Z�Lw�I_�*��76f�;�:�a��(�zy[��#T�g��~�v���h,��S�V��{ԇ�N>�7Շf���wG�Z�r��_cl��,CD�#��	�F���5���(\|v0o$�#aw�bq �.��!ɛ���tw�O���m0���E���������ޙ�gާtG���+V��EŖ�rӲ
��ތ����:��=5���d�nS��&]5�V���j�=�9p�[�-�� ��vg�x�4���ڷ�@iK	}�߱x��d/�#�3��ʄ�l���"�C��Go��JKJJ6����4�s�5������XT�����bZ,RŜ��=u���+��G>�~ASfC� Z��ԔU���8�9�~�T`+�Z�B��L����RP�ڕ�J{��N3�e<0bG�ӧ}��̒փ�'���"�B1k��Տ���#����&�<5�q~}z�e�0s^w��������&ؖs)g�;*��3�g��3��M�}];�ӳ)h�䞨N���>ڻ�%,bn�pB�"�Bސ͈�ğ����tv�ff%�)*�g%[�m_�#D�M���i�Spnɽ0/zc1�j8y�XV	O�X|�<RͰ��v0�(s�+��C���5�n������ӛb���%�ҵGN����s��@`��-�0l���ƭ�%R*����g�t�C��D&����m�>�e��צ�2�&6u��W��O��.�4|���qd���>�6�~7��\�S�3����Z�"�����|���ۧJ��hv穔<�1�?o��$�:�ڹ����4
�x���7G��i&��g��ݛtɮϖ=��=E�;���05��@6�K�E���RD�q6۲c� ��Y:���R�w�?���t����8k׭=y���᣷#�������G�f�R�j~���H���HM�R{�ܾ�,}�cǜ��c��}-�iv�q����ܻD���u��n=��uqo�^���)~vN(�b.-w��rI+��Wzߑ���3�x���k
��͢u.��!��^v�ҥK��@����ގ����T��}=�I�#�;'F}j~����?��y7(�m�ל��_k71���/l!���wH�]��լ�<=���	�GT���~���#G�d	)e�nDRb�z��j�H�w?�.�l�I���l?��m�[���I�=Rк�"�F&3�u\Nh ���'`�U�/0ia�����h�mi�#�z=�K7�6h�r�$ׇy��uh {�}�gdZ��^fg|f������L��������Sͭ�v�I���p�Z{����vC@�O�vdXrqH �ؒN
`:���5�96ԉ����2�ҮN��]688(Dּ�{<W~mSW�3׶ Ǐ`�߷MeΦk�EM|��l�ӧ�rH���A�lܴi��yĊT8>3���m-j*�N�4�yl#_Tn0�_KQѺ1����X�#a�h��5)j+��{�Њ����8��B�����QP��{��ro�����0���x�&�N%���,�	mN�8�m77�Y.�a����/7�>���Y�V��^�#�[,�}PpT��6��;�?�U��6��bY3{?b��o�Y�(�����Wi @�q�Y�,��m83p�þ\���^z�;D.e��*��rX{��ޞ�qg�����}��:�~\ץ�w�����-�)�-|uv�[@��\z\��=L&��N�Љ��p�`L�m�1���g�,��mrt��og�8�,G�v�C��ԏ����P�:�d�J���ه��0m+�z}�]E&��@8��-a�������W�tF�k�񖜣�v����g�� * Cq��h�#Ge�^��-��Ϯ!+=��P�U`P�<� P��y��-���v��(V-H&9��xl�Uԉ]]ghf����.h�;w<�`oГ-&��q���I���n�n����壷�{����	.y:M�}�����mHWϞ=7�i���P�Fi%7w�2��7&/î8�h�<�S~9�)���q׮]�N~��=����WWz����b:�~�:~�*t���ם&���2X0M1|��X�x����L�r]�&�Ӣf���˗V-��o�s~���Gh|�nP[���S�� #�U�uNՂ��ګ*F��N�w�0O����s39��,ԙ����\���^�=o��YM�`��d��:��w���#��i ��Ig%�=�+�	L�՘:�@ϔwd�ݧ�����:��E��&}D��':����6�17�-U��)�5ܰ�w��=�Ik��:�+��}����������4��֮mAR�^Г����:+��ڈsv�7�lG5���s8��ҲG�G x������CJ�1�I{�-�;2#^4V�j���B��%�nKV+������~P���W�ק[-�T�Y���wc�}̫+�L�Xԏޞ�����N�r=��{�����{�b��6�Ӌ�a��:0��G���.�B���엫�B�Adk4yӬ�/.d_>1=� ��Zq��/s���O��TVL��	!�pPf�h���]����v��7r���P�tn�ZH8�k����w[�;+�u��-�6+@�uD@!�G�*��[�K�>���T<�#D�q���'�g�߾{��,�\K��ಮ�.��x5�u���ޚS�cgA� 3ܴ�|E���8rğ����>7�����0'���m}zĴY�RG��=!�i2��Q��I��;.��M���z���ɲ.{kRN[Ը?�wf�]$t��:�� �����vefL̄)��~�4�Kwdl;Ƣ����(�s�:��
�6L8��?��q�Omm��sC��,��w�c{�/$ކ_5��ޖ�)5pq(��rF[�b�<�!D�!*��fE��A0+�E�����ή��0+��5���ka~h��bX�������e�`��l��+?do�9(QQ��n�����q�Ӟ��ys�9�6|2!�k[����)s�ɷ��S�n��W���]��OI�yl���M��ʙ����e�v�M����v�����y"�o�)о�J`z�~�+��E�ne�k�Lм�)�v�����b��3?��3��"ϝ�3n޼iL�^/ϦF�[�j��"sh�>���.����wM�\z?:2�����~k��&Єג;�������	���8P�������i�b�6O�^{{�� ��S.����ۧ���N,�?��i��D��4���v��?ƺ�٥sz?0j�-���r�~�����]�~wO��~k��|u�y*���>m�zfkZU_9m}_�z�ӟ\S#���}�L�uS`��C��K����t
�O���+'>8�[}��B����}4�F���^�c09�EN�ܪ|ߖ�{䕹��.u�G���I���{��3�%6�w�Kk9�T���^_���������{:��������^<=|�4]���ze��iͥŮ�5�K��ܖ+����~��݋�A��N�;'��ʾ�ǖoy�k��)qB���S�
~\�H#�_�n���}3�No�������}U�+-qu᪟u���]�����c��9���e��ү���z]I?W^���d�9`�;�H��v��f`�ڟ���J���?�_�SjYn)�(OW?�uN	M PK   ���XP��/�  ǽ  /   images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.png\�T����"  "%�R"��%�]�J7�ҝRҭtww�tI���<��]wݽ�Y.����;o<����U�GA�C���A��Q���u��y���s}X��y�($����������H����,{;)�z0�VP,~gN��,khm�l*S�6f��}D!3ܤ��VR�q{�Y\ÑV�]'A���fӵ4�ϓ��q�K����y���q�=~<I�����ӗ!hG{��%�M?�ă���w-&O���;z+8��Q���f���~O�&��D���?��e�yJ�@�-B�����z%1�����>&]���b��bp��W�	�H(a�o��d��-���Q�+4�R\�xWe���*.4�����oq�`��F8��c�L{p��ڢ��}
sR��z�S�!�����w�
^~&�*]��R�\H��sݐq�g�A�*�{��p���_���tcd�=㬖T[`��e�b�^Y0>Y��҆�R�L���y��up������$:�+􇇇�q2o��h�ۮ|�6 +ݐ����%T��0+�U����"���7��\��A����'��KF�R���������Jy ��a��υ�;�f��J;��	}|��j�b�i�]�|$1�\��s� i��~b�ͤ=,
�Ȁ��I>��[$�m��-"�c�V��g�~���'�����K��k>:,��.�"C����H��3�_$2^.<�U��)�	W����
ٟ?���*ȥI��+̕b����b�
�Tm&��J�](H��7{���w�xc��%"ҽ�Q�Ύ���<���Ͳ��kNtttfף%���qj�ES���.���8��a���A�Oԧ	�XH�?�����K���s� ȸ4w0��.��\�g�?��涉�Ȃ�E�L��/ڿ�q��1�w�0��ßj0�������@*����8�����E{gm�R���AY%ߣ���<,�QO}�o���04��=����_/��W��"BB�N�l��0�\@0~�h�U&H$�=��?�W��� u���YLAL$��Sh�,�٩�ha4b>�<P%oɁ�@����S����ez�R��M�/6��C�i.f�����oӳ�������S�ae*���r�|%�|%�MV��0"u�T����B�l���2w�$����u?I.�ꟆU�nn80�����00x��0�������CnbȚ	3y�6��7P�_,��
D*��{y��?�%���&PRVN�!��d-O��6�_d�����ѫD��,��V��c�݃�k˩�$^����96�
Ll_Q��z���)�����%��'.�7�ٓ����>�$g�_�1vm����
	B�^��z�t	
��;"$��UU����.���f�B�փ.��'�����뙓 �vHOW��3� ��S/
�����?vW7��KF<jF��Z�G��p�����V��GF�;�uu-7K�Ɉ�(!�a]�"���T�OM��<7�DE�待6���V�!�iJ�%9�f��f�����S�?2ޤ��CNS��m��^�?=�b��vjwZe����R>(���/�%�SF�'�g��a��渶�0n�C6�l���_����o���ͽX"%ُ�
����cka��,x�|t�|rE)Q���;��Ի�I��_[���W1Նp���eK�w5���b��k!0TW;O�/:"��M���{c�;�_�|E$��E���+�eE���K�k6��	+7�-��I�t�S
�^�r#^���Hw�k�����!��#�#�k�K%%�<\����D-���M�=	�F�dq�8�455[|�$��42�˖�p���c�٢Q��X^E��\�:��祺���Ĩ�sh��7n���sj���i(2T�E*aY���;�����LoD�Ă��G�����=S'owk���K-x_����>I�����D���Z���Ͽj9��!CO�7���{�K���dvu�o�W��aA�sbaqS)�1K�"�w�Q�ӳ���,}9*�΀���4[(���8��`��}�慀!.�?�XT==��0�*T6Ư�"�ڃΏ[���l%E�R'fH�p���E�� 4a������ײ�|�b1�c����aID��9wf��X��Ku�0���d�0��,^�c?_*��+l"�.�������k���Թ����ܽG
u.6%��M���
br��O$�N�?�?�bi���ܛ�\~�u1t`�0�AS=���~��3��e>z�����������uR�@�h�|Y�+�9�qM47��B���F8��&��O���\�p�}����uJ�y�H�k82z��_��9�"�5��`-��|&r�LS�Q��+%BŠrV,*����#om�.ל� W,�}9�@�p�H�����'����P�6�"z�6���?����aF#3��|8��?N�~{��;6��K���14��p��% ���8[r��N�Ȧ�B/��W)���e��ckm����"6I��ߺhwFDD�WEB��(qM$2)�X��E�/��$j?0T:9�TU��0�||��M��sC����(e����jZxU׷Q�
�}��i����D�۩a�� p��	�SvG�'<��ƾ�ãV����	MM︤е��Xp>��%G���*ӕo�"]�b���Õ�P��el�{Ԙ�� @2}�HI�X֦����ݱ11~7�;w�����YR���q�����&�����hn��,��Fg�؇V�S�^���>��.���4�榤}��������Ot�"+~j����"�%�`����W�
}m�?eT���u͝�_�Z&L�F��CDL�����9A*pkkˏq�pq�⡮���?�xW�I�v�SR�S:���J R�U��0�-�u�T��!c\�W@;Gj�p�Ic�tdd^��6��H?�v���_c����Q�C�� _��\mh�,,ts=��D=�T��_��+���_+��1��"�.5Vѩ�0�9�HW�
������NŰiL]��㝳��ԓ߆T�b-N4�X�!�ѥ�*7 N8h��׹��:���0�OOˤ�_EtَD�b��ţ|b'�
ޞ���QȐc�7�bq�b2_Ǡ1Nhc�1Kp�,�P�Ģ���o���F��� R��r�eU���mWa���Ƨ"�9��+k��uZ$�*6�Ud��Y�̪�a���W��b���K���t�<iק�)Y2�p����Z{[l���;=R�Kţ;|6��x�Â>��&�h��L]Q��ȒQ��W��\�E�����8>�A�����,`�E�� �y��7����YQ,�˧6&~qk/^���m�(�M�X��O������_�.s�E��L�n��PBv�l#����c��J�&�<������,������>ߧY%t���T�>�K������&t9
��چnA;���	����"����?]p+��hm!]��r�?_I@9u��g
G��\#��Z:O��0����5V?_|H��
v�x�&j�\ϥ�W~��s���z�ֻ�!����	Ve[�Su��梦���{����z��l���kr�V���s:����G�M,�<t����ю�a<`%
�g8�/�lG���'���n��.���y�y�0@�Ȇ|A��[���_cbR��"�pj�;�=iD��YN�Uv�����a|?<��1�+���ĥCA-�c�ig������D�DDV1�-���DMArѿ�_�m*���������²1X�M����X�t_����05��0~Ã��<��m�=;�M|�1y���ъ��݇fB���f�R%�Ye��4�i�S#�I�{�y��{���ȗw�#3U��~�#&���ԉ�ls�S�����Jb!v�Ϋڨd�{|��a��b<���0
��o���ajb������n��
K��gr8_f��/<��W|���V��20�"O5�T!6i[m��Yk|�Jhy���H!x�%�A1|*�v�C���h�h|j޿U>��Z���'��[��v+�bnv��@S����Q.J|<Mn�";�o��Y�|�[�o�h&ȩU��Tc�p,p�Z��ҼS9|�B�e�:=S�e�o^|�Or:;;v��I^��K�5^����.�͐�ު`�p����E>�á	E^�a���0~7�A}�e5�����.��\�dHu�3����ol��b����1tl��I��?��ҿc�ś�BQ�1(����"Y(��W�����=�z���7�Y��mN_5{�z�,
&�������9�\��і���-1$�ez�M�o���E��{�֎Kߞ��b��s$�J4�v�?=ɀ�N�:���Ԋh�J����Ս>N)�CJ�FW�%���iq�t�0/Z����0��X_b�ǂ��4����S��J(DG1ĭz��.-��ѧk�qpK(1Q����q�]X	�"�C��vf���*�Dy�`�����ǳ�!�-ň���C�/oq`��Ia��f�K��4�s�:�^7a:"���\�+{g���j�G�3z��A��+?������h��M(C��v��[�NP-&���{�e��O���q�!�9���>��>4�WX	*I7�;��݆���V�5��� H�*N��zB�I��}�Z��*�n�ӣ^fk��22�;�iqf���O�n�%����$B_&��W�������V>���o�Ҡb�W�&Xߙ6+I�RM(w�(A�`'}7���t+�sC;���x�������.S7R����eQ��f�&('�
�� J�&����FM
< ����U,|Θ�JM�_;�p;�;���N_�^T֩K�b�{AU��6�1�.5W|�����|��WX?��՗�|�N��y�lyk�V�����w���H�&��W����VS6C�+_F�}���5�ɪ>m'�Uźi��9X:(rJ)�����w?��Qu��!>T6�.�DsTr.jvt�|���k�C����\���r��~v����.�B�� �G�i�xJG��˗<3�vv�F�A�B賜a"Ga�_��ε4c��ɽ�:6�W�M�˵��B9�q������~=M�n��8�a���������[�P��
���uh�����A���g��vF��zk�/[��aM�������L�sR�ӏ�Rԯf�T0wE�3�Ԣ'�jl�;�0ˊ�=�6�3AuH��������0�7��F���XKX|E9#).'��FK��
װ}S���nǂ��,��jo`�Q��l+*�f�N��ox��x<U�����Y'��2�P��sɄ*��]SַHf�t_�!ى"B+ђ� t*� ����W������7p�_K�UU��Ⱦ;
�<MWZ�1�r�'���$��R�E����1D�C=�Yi1����U���_nC���	�d޲��?�h���:6�QJ8�vB`Y�CjP'8�̋���%�D<��2	������:V�`��<�#�<��P<uK!�$�Ԍ-��ѫ��@>@�v:��Z��n���a�̆ONl�_|��Ϭe�2��BX2Spn	z8H�P:��r��N@C/V;�R��9-S���|�W����*	�m���
��9���!�^<E��#9�%�!�qn�Ÿ6&�4zU]7K�yQ0��ͱ��?n}^�WW3O,�K���7&"�S�#�>�«���p6�LN���/�2Ďywtq���$x���S�������zh���@�ʾ��Ef�S�Wt��z�e�A䳴h��F��*���a�)(��
�
�mT&��M�o왧8������n�Aɍ8{M�6�Y[�u�Oq�ᵃ�A�׌�ڴ��RMK�-I��m���ϘõdT[��SW����t���*N�-�ҋϲ;��%	ג741[�y��h�"N�,�_P󣄗�V`:��hS�xQ����j�k9��3bCHԓ�{Oi��#{��dm�O��	N�<�m59զb��#"����ܵ�q�[g�x>�M66��ZC�h6��?]�K�X��c��ta�p4{Le1e�i3�<�~�8{���g�,
"H��Z-[��+*�3\��1���~/�s��K��Z�#qܢ��&�����~����,tO��
�0cبu/�(�U9��Y����Z8���һGBԭ�g�v`��$M 	/Ơ�2�K������N�ևr�ބ�1�ī�,�k6��g�^������c��%x�//EX�{!h��t����;
01��,P�<����.p/|� g�t��q�)���od��em_Y�'�3l?�熍���4�pm&cĘ!N��3G�ێ�����s�j�3�47���~�B`Ts�b,ω��-����s|l-��r���X�غ7:�G!#��n.y�8���)wSj��C�_�*{�1Jʟ��Nn83�sԼzы�ɕ��F��Z^���K��Q}�i�[  �l�$/m��D)�HH�YZ8�}��]~3�=�"
=@�q�����L2e��PF&�cr9q<ҋ��d���-T���O�����)Y��0a�g�ܟs}ρj��`�!&�mX~��u}s�"�M��n��#ꀺ*���}y������s��I�>%J���d�_#�=�a%oV5������>�P(�ph�˙?��K�rVm�/�Q�g�2?�e��gɏ
���xk��f�N~]�����hE��2*:XF))9#��p���bz�3�|�~Z����16���`uLL�_�����}��H��^���L�}��/�!Oo�?�Z���n�����kG�_qW�}�V|��y^]���t��Q֍A ��領>{I�P�c�&�"r��,�R�S�{�=^��?^��q��[fy?���k\���r�|��F�]�ߘ֤S�_z�6�h��5���S�v�qYzM��o�5��}k�noǙ���Y<�C�ƕ����/;�r�T���Զ������\9�9����}nH9^y�O{=à�'e G��|s�iɴ����M��f�_�X���a��m����r!.d��C£a�[x�Pռn���[�b<���L{���Oq�U�:��Lz��F�U�9�$�:�m��#��M���Q���޸Oدm��>n���[j��Q����k�f���6cbZ9�}CU�:�s�vpJ ������s���oƄ+=y���W�%Za��<Z��ڹ�/2Ƒ�K=�^�������gJ�V���A��v�����K�#�ߦP�Pf���p#U��.2�ϛ%n�TsNy�v��~ͯ�w��=�f[�p�<���>S�١s�|	I�&ˡ�P�	�[�\u$5��1߫�;5�������}��;�l� ���S�jGؙEzI���F��2M��s�7�9�/�d�BBr"bƞD�A�Tn�V� �}��t����s�)�
r���K���F�����H��hDov$ټ�,]l��>�9�+۠����z}�n�H�ȋ
��ʈ-j�"���qAl'��%gA0�ϸ���_���K�tt�_;K�*ѣ0�dh�2X�ęs�n#܉|/7�@ =
��
&��G�t^��:������Pa.&s�:F%!]�m;��pc�[G�'&�\�`���J�B�X[ִ�7ϲ�^�H��+}l��U���;\��rg�w2��[<�b�;jo���=ryCg�-���d;�q����)�|V-8hޥ�C�,�XVXH�zG��I�.k�4��{��Cw��IG�篫qK$�RT���oȴ��%X�u�2�BE�#!R���k�J\{@��p�	����(��j�9�|���G����Ifz���V�곾��ϒ:�Z5��n���V�܏]�ֵ�_�a�����lN�f+�d)�����(�o����C�;��Ȭ�0���k�	��_:&�lcH��ly��:�~Cn0�޶H
���\L ǁ���b( vlG-�w��,�������_�<�����m2�;���}�#C�v?���9�K;6od�mH"ÅV_	[��A�|��l��'iD|&mn>S��j޺�����A@��M-ox��v2��߭0���v	���� Z�՜7�dnP�7�|r\
e���f�F���I�>�Ev"Z�$�e��9�O�8^[c@0��0�UU�l򎸟�"����������酕ge�/�Xj�q�N����X=;#�����rP9s��=
��~F�U���q�dd��Ё��o�����v����ԠayRjU�[X,Q�D@�O�Bd�=��l�fF��u#�� 6O)��%���_c+4�-�E>qڋm�������8� <Hd�߼ϕ�Q."q� P�s�pG�	�#̇�wq�x,�Oi0Ϻ��7Bf|ۺ����*Z��+�eQU�";[�=���f;�3���-< �E���p����( Ԋ�E��J�]����ec]�B&�++6D�d@n�p�ĄH�V/����9`m��˕�F������hkk�벽@���<�
ݢ���aT�0.a~���V�"����E��iPnp	�ǭ��beU��+���ddH/��I���?K��N⯢I����DU�eR,*���8(�H�j�

&���~�c���՜��7s-^,3[��6[s7�h�,h�5J�9��
���k�*N�����3�P��)��C��`�nYD������w�CZG��jk3�j�������{Wb�4��`I����B�Vz��i�����5����G�D�t1J���$�f�5w���M|v08:|�����t�7��p�A�R'�h�d�B���(AG	����-��-\�FA�b��j@BԵ	
4�˝�V"x`kB��]��>)��;A���0��A߶DZ��t�@C@i�C�_�*��mmS離��i*��-���qI��NS��Qx�����>�TIB4EC%q
��=r]>&j��Oh<�u)c3V�lb5�S4#:~Q���}�F%���R��u�DQfG�Ǻ�B�<�c��	�1��^|�r�v�X��w�3*��V�����BPN��<fY��=d���U���S�1��t�K��� �Q�l��J����h-%�CWH�~!�*n��v̞��ݶ���MP�ٓ���h�i��]�����Mg�ITÈ1#XX|v���j��lE�r���,L�Y����6���v�g�������D��bK���J\�M3���q�H�~a��Rx߾$�3Z��Pm�slӂ�O x��G#����u���A�L�����F �C 0�*����� �]�.ߋ���E�E�:]e���R���y{�2��Όߓ��x._�z�At�f�|������'��!��/�%4<����-S��A%��冽y�R@�d�rL��5��E��BlR`	�|��5R�^�7��l�1�w)Ӡb}�0���GD�}ng �Ɣnӧi�F�l��H<��j�R d��$R0�?)t�1�=O���7^�╍�2k"��џ<�L�ݿ�Mk.o\�Y[.��jY*������a�M�M2ׅ�$�~!�	���0�Gy����]�br%/�|��^;��(�� &^�<��1��p����Z4�`��F6�T7�k��G#��p"�D QFz��j[�z7�G��n�cpS\� ����&^� ���aM��k�D��v*V�@�mù�("	k���BS���od���q_?��9획����OP�B�I��+rY�(�l�:�����zL�"O3�*����qZ|��u�/f=��`�b��@æ� #q�]k�?a�)~�򶱄�h0j՝gǮ�#vIdShIs,���˗����A�PDz$�~�%�����p�-�C��G�����w~Hbn"+G"$�w���_k ��[d˻�����a`l�����_!�����Gf~0�/g��[���	AT(�jú�(�U�l��g4��ul���+��^y]֑ex5��nLpǐ \"�.���u�RYLA�, T�3.݆��Z�q5(F>(���:�|@��ٵ��}��[���LN���
�g���	hh�ҳ��t(�T�HI�)9Wq�����ק��IP����V��ܡ!!���!:,�1�	�B�zj6�^ ��c���I4��x��$�4���O�k��JG���@ރ���>�K���ӈʅ��B;u��{
/����S2���B/���{��	_n���}�����
�d�T��ٳ��?4�@a���]��*�(������O���T�ȑ��`�HU\=yr��Z�X��an��CdD΂�����4��5�#J�5C����D�48I�]r�n��r�x,�
u �4�w4x��"�X��S��*m4W8- ��$��+����}^�.}���"��l��S�M��pP�N���H��+�B�VbKq��������Ҕ������n�.��R�b��V2@G��=~�a �\-�BA���b0��>��� 1���5����A�����sC1��� �D�;�7_ r?m�4��~����7H}fx
���~��Z���~M��9��.�*�nk�x �5;�&�y��*����+�`�T����K.��oD��x�7$�ut`==á�b��R����t6P��Ǐ�B����q��]��'_k�R^����1Mz��z��Qf)��E"����4��C0C�>�<��yE!���rK`Y*�=�$^����T6�Xɗ;�%�JA[Ԩ�[mH�m��Ph"�-�$ݗ<�pt�)H=)=:�d𨎿N
1��߯ 0�Ej��\�팷q�q����s��p��.�~�b�y`Aa[4�J������"Te�CP�����"�9~���=��g��9Y��B��[&��Π����e�o�����-�3���ǳǾ�h�UE���9�
�ʐis�Z)�#�-h�W�� '��]2D���&���Gƪ %�02sr$��(i�d\�
�1ެ5����(���X���ڟ$���T�li���X
�R ��"�o�l�FrPQ��m>\�MW����l�cn��e6YT����_I��8�����ⴊ�:���)t�tj��"2�J�ۗ�ǃ���������Hl�K+~@΃�Wh}�Wa�<�4 ۿ�ݲ�3i�"�C'*�DT�^i.ܱvۯ���>�0�B ���z����=��:C嗣&�&>��C$iy��>�<#;x�vwե����@�]x��#���<孷���j�x������f� zX�S�aB�&u �z�!�V*�$ UO��b�X�Vf/�l���%�alBF����騜U��gi���>4�kjj��Q~92�ߒ���HT2�e�.�X����# J�s��y�l@�4�. ��4k�&��>hd:� ��6H��e����h&��c�T��b�9��t;#{���#��y^J$n�h���z����J�uȍ_ݠL[k5�e��qH&zn/����A�|�����������<��a>�ջ�l�f�}��py�.l���R���j����_8XW>!?��$��i����s�)Զ�u�+o����6 N	�s���ɀNl����l�jP�K3��Zt�TPnj��g��9G덊@e�(x��[2-�HY�9�Q:�I瘠��:1ǫ]�G��0T1�T�z+��zf�鿻�4��٫8��K�~`�F
F/�0!"g��D�����}�5��Kr���3X��	�2��uv�趆��S9��A��Q��Ȅb�L'l�d���~�]Ҽ�t3�~��O���.�>H���>9�Z�j���l���c��l���؛zq3�O����f��o�cي(+�~��gVB��2�K�)\d~�HHA���|�T�%^
0g`G�Ĵ�C,��B����[d��e��w����w��7���1mh�2��f(���Y��m��xs$����9�lr2��-��!f�!7 l��I����N
D�ٽl�7�K�Φ������oV��� �<�.�*@0�{��i�E�����\K�meߗJ����]��.	������?RPHHIHII�ʯu=D�XMՇ��ݑ���A;a��!�ZG����%Wi*�;/l_֐R԰7 *$OE1O�A� 3�&@M�
{�G4sds�]�a�VE���
������l��� �>�Oh��eyPJ]��]��Q[]�,��o��b��v��<:e�-W�Fɚ]��[�a�Ҹ9[� ֪�=��Oz4#�l�lRX0�K�1� ��z,�4ğr� h�V��� ۏ�"�-��v7)�Y��zRH>`+~�wfO��A��#*_|�7��wbc�I%�"�h^`5Qv�{�б�����8�e}����׸#h�/:����t냆�ҲI(p���k'�&�^-���H��<��}o'��S�t˟tuu-I�ɽ�ɋ�P��@��v<C�b���8�j��d���ː���w�j�4��ٿ�L�I���m0$;W/�1�@
A�V�p>2<,��H+<-�Gl��hM�'�f�)��b��N���#4m���8����B|���K&��t�8�"� 9�L}� =�i����+�b4���\*߫�]̙;������h�ɐic� f���\H���0~#���:��[Da�9�hSq(�Ua1��R����1����M}��@�5g�&� ��m���'<���rn���oR�#��6RZ�룠9�!Sex�p�C�[hwh��UX85'&���'?�����$���:x��vҐ݆�mG��o�H�|E���"��X��~��l�``�@S�����h�X��΀K�$Z��s�X@���U�H��br�����E0/!H �`h�3���a�ێ��O�j(�P��%6O��IE����J�� �0�p�n��u&�Ā���*�}
H��_ł+!�m��݀��*�c�@�+�7�����l��X6˭<�;M��$�n;�e�x�Z��g���ԧ��Il�+�F�m]rh�� 4C@AF����a��6~8
�#`f@�7�)\0���4���<�P �$��X狈^��a��� ;��n�"�l���-�yy��G�dn��� �-)�~�r�x� ^��?ˬ�a�i ��Ѐ���L�138����4�����j�Ρy�l�h^��������	�J��6��Hb��!���`F��i����W�7E(��Rm>��� ���^d9�p(wt䙙~�LGճ�d���	A��ܮ�꽏�����{�;mp�6l�R�1���2��_{e�Jv���(���{ ,�U���!����)�X!��ܚ�(;�~�2!
�����Iyq�E��ݍX�A���C�sw��\T�d����~���9����5�)�l`��90����כMX��[���r����"�#ض̆��r{:����^��z8��Z]�r>��|�
���J��z���ɝ�H���������_�X�x�p���>V�3q�S�WP�T��S�����v����L��f���wu.��V�{�v� a��������g�L���gVi{��,�X����9]K1v�����κ��l,���:��.ju��d��&�Ϟ,2���]!���i�.R�U�i�B;�mFf`�+񽮸ѝ�u��q���Fh�c1N�n�Ϲ|;?���b�i�n}�	���,c����<��O�$��|�5�ި:86. K��I\Q6�yc	��o�r�(hIƅ��A���W�����}}�㥠=.���������m�M�
?���;?^��U�G�~QR�����Ix��	�[���+�_c���8!p�9����y_����cp�j}��p�PU��if������4}�������y\-X~���Q���@�ɝ���+���_j-���#�.R�о�[mkݶ���P����G߉cU�dBǎ�����t~*�_ʨ����o9��M�� �g��r�w���5S�xd�M�����C�zǫ�A��k[��w�H�Fļ�h�Iv2�^�U�+�Ľ����^��00���k�׉)z�F�UI��F�=Ӷ�׍hw�=���\��5dw�v����Q,���r�����;)���� ���2���i[�E{�|;�5^�����9�)�U�-��}&ZS��k�z��樿U^�~�dp�d�r4��u{CJĞ���v��nG����K�����:���@�s�{G7�:���v����ކTW[+�����Qu�[t�I�jG�s>�X�ٮ��8�hEn�~�pGl}Y�_�T<�{�~��\{Y�N�&{�� ����dx���Hq|��w�_�mџW�OZ��%�=y/%�;����W]t:���ӕR�ΰL|�'��P���r#�-F����5u��7Ew{A����˖�� ��yΆ蔲�k�b��}�xû�����Ҏ)��\s�q������ֻ�ޮ}7������:��'Qt�V�7�9WB�O��W��s�.��Km4j����lfD=�MR�6j_��16�-���[�v��7�ٵ&>1U.{��T��AY��u��ߛ�%�h3j+�������'%2��:��X����kk�����KB�2�}s�f���������'k셣k�4q?�8���J�l�%����*4���6��aN���6�P��<wĮ�� *����*7`��$,u~�p�&��=���B��/�;"}򑢵����*=�{�|ԅg#�Ѱ��-���%�$�H<ߓ9!�fd߳.ץ�Y�fd�W�$s{J��AM&	pG>>4W��p��k�DG�l"nsE�8����f�M���3È�' ::����!�zafn!p U.�������f
�=, �+y�e*zW�g zqc4`!O�Gs{��67G����z�&-��r^J���+�$ex݃� 6�_��;�|�}|��wW5p���?�;��+\Q�h��K��L�N�|��滸�5��`!�޾ߴ���d����l�8�V�{����W,�]]��u�����(*	Z�o��NQ�9�/�g��6S�ÌA ;�fM��3$`W��\=XhQ1B��m{�=�:���$z_\i�{k�E-�N�ɣ�����,��:������L����*��E��;׾Q	�� ��(�8(�G<RXI-�S��ߒ�6����4�\��j��|����CL%1�,i��J�sP7	����>�i���R��K����ۻ�M�)�g��p�ܟ$����~�/���z�Fݥ��HV�Cj1@
�]d����V�W�I��l�X�
)�np��\�l�˩��oT�aaV�����	9���Ȣ�~����`9�Ǧ#�M�Ǯ��.BYu����������cH^ �74�g ��eEFwzb��7\R������W �$-��κ�D L���%b��	5���n�&�[Z;)�$1 	��3A".�[?��
s�^;��/�Y�@x�VR�����0;��/CO����1R��
�Sw��8|U?�b��g�O�-!n�p����灒£�?����5��fx��4y�g�Z~��yU��`n���=��x�>��¦�*5M_6�﷿�o�uO8u��OuE5樜>b�94���+�n8c���+R{��|�V~N��j	9~�on��ڃ���ѝ��Jg��(�%����]U��yGc�[9`s^nJ���'	Ԝ��6�t8�Z�ޓN{��6����,*~
�̸�zƛ���P�H.`Dt�vBD��^��DI���S���-O��PVڽ`k���Y��C��Ư#��w��ʮ�u�,�P�jGy��ߏ}��ke�O~�捎�6�5�)�֢����zG���֚�����B�r�"XQ�o��uɅ1fXo��PX]�[��7l��pY��6�I��w�i�z������v��J�%婻oa�E�=]�.�~�G�r�?zJ��4r�H���i�00N���#�,Q#·^n2����6���8 �$B�@�L�}�b�^W��(��}~��dZ���s��Ni"��Od��I����%�8���/O��/糿���?�sK�~w/a�e6��U.�"
���n�ϒ�hh�b�a??�\���h�Q,zG�S��`j���)�~��
Z�y��fѺ+����#ꆸ5�ݤ"������sLWy�������qP'3�T�F䥝����(�4��X�~��l���ğ��t�,�V������]�����W��G�85M�.�F⟠�heU��p��}WUK�?�ե������P�U_[ˌ�v���.b�+n)�n��<�]��?I��$�@�V����uճ�(�?~7��L��uX<�p��7�N3k15Wk�[��Ѿ�k��j}��Z;n�h�?�н��8�e#���+*ԏ���Y��/��N,ե��ȼՈKm�G2KҎ��������3Α��?��SRo x�j&��Y�������1�����\9I������Z����:LPЂ���"�>U���	�*�����O���'�ӛe�y��}�Km���gEX<H�w<n�8c4�eE�H��������M���XZ^�֖���=�3��P�� |��������NI����ZoT�G]��kn�6�t�ܑ�Y�����g7=��^!�늀T��Oq�s�B����$��l��c���/����,R���ѼՓ�]����>��3��(�[a��@܎�/����N	�3�}� -^�h�x~�� �Q	��X�%�/)�D���ao��S����o�y+`p����8��Z�΄]�ُ�؀�:�%���6�.@S7��G��H��.Ȍ���<@�J��e�A�>h�#�'�7�;�ǫ~�<���+Ϭ
_\W�~ݬ����'�~ʓ���l� @dx�uk莑�9=�]�v=sH�����m�ĺ�%�\����4w�Oy����g]xz��48��`�[�nI9��z
,��׮�]{�h��l����o���v�����޿�~�ޘ>�^�Mx��i����W%��ȍ~����p��)���%Ĩda�'rh10-M:6i�� cfA�)%5���>� �y _/ ބ��N�o�1�r�dg�o�|V��5"�ܗ��]�k$y�2Y�Ji>�#��A�.6�H���_�]ND�H�~&����@���@X�����T���c6��fܴ�R����\�)�C�l����z�=��QT�\��V_�x�죵����i�\��.�,�f�ڽ���2��"0����&�Um����T�OdL�S��dmMU�Q19��(�c Y�<����<��p��w;��C������bzV����|6z��Z�0H�AW!E,�8O��Q�F����Qƪ�&,P9��9ƠkA5���rG���W�f�r��y�jp*��~�%��CLP��A����|w�����^��+d�C�~�	?%��d���+e�2�I�����o'VL�U�M��W�?��d�]�{�1K�i��J�~8��sᚳ��s����N����h��{�ㇵ�������{�QA%DDZAJ��K��E��`�!DA��`讁�������{b�O�/��Ď{_�u_�ޏ�E�WD��Rx#v�n~�w�I��)��tR�m�}��xFj�tߴz���,�%.�[�@1>�.4~�-��]�g�uY�d��؁���|BYfB��?�,G��{Kf��d��IG6���(g}����"Sީ�t��eyGz��]]�^�~.[AAM�I)g��@k@zԥD�MQ��L��b���c�D�`_w6�U�f�����9�޹�ܪuW�}���4S�"�L#��J�#!Y���r��;>O:���E�%=��i.k���=m�@�1�ː��:46T�@sQNoma�^�M֔��i=�a,��;h�AY�8��M��@��pM�������C@R�j�>qZ�j�$�i�����<h���1x��L�pM�/���?��K�(�^^��T��r~18��~� ��#�HƵm+��F�: #ؑ��0Q�6�P��)���W)&l�_MT��,�0!`kG��^�������w�����i:��,Y�]���D�(�m���I1f�K���|!��"�e��ȝ�	'�WǵU
�r�ɶCЧ�z����@2d�3���BuV�n�}.����]�1T���8Ʃ&k�>���Ī0I���ًY�l���9���wQ�K˔=��-�x[0�6��#w�����KX���_T�f�S���i��#����_�x���(������O�~e���<������7!S�xSd���B]���B�l;/[A�;oWۨ�t��ݢ�����[ߚ7���9>��24$���G��O=��D"�Yyޛ�2kui��b�׶c��?��Iې��yr&��&uT</ ��"�o����7�}.'�j_W;��H�1ez�E�)fd�E��	�͋�)~@'�ǫ���z�Nļ�!j<��"�@�����۩Ǜ�i<[��_�}�J渗��-+��g�"�Q�vIVWF������C����a����W̢�Z�|�&#�p���X���rb�˚�=Å���e�	��'�Q,L;�[�2�_uE>,����}�=�Lg
6yx$��4�$�5k�A�8�|���]����&�,]�c�u�w>����.�~�ъzM��bi¹[��R���d|×'��(ݽ=��䡯�b�����7N�)~�I�$_<�rW�u��划ĸ8��Tt/w%^��N���A��bs�?}�"�	x`�ř ȍ�W�����&yDh�_��:n�����?����2�`��Rx���-G�S�Ǩ�L@�Ȅ��i���p���S��@��j��Fz���Ț�r�P��;��|�w6ў�r�NxkBN<�Z�NtP���$�jvH>�����~���`<!���ne���ځ����@�����]�:!B�1����!�s�m�Y���r���È���mZ�Z_�p}t�ޛ�f���9��"�Ғ\:�$O��pg�>v����k9/��B���E�k��Ne ��(�`v�E�$wt��f^�]=U�Ć�Q�S��g��F�ٳ�y0��ލ���h��1n�
��N��(E���<��7~$����b���g_O/f�N]q�hH[���M̆�# ���� Ͽ���]��>/���%����EAF_����)e&wa]hI|h��eߛ���gKk�J�mׅ'������ќ�%�PO1��g�@��2�J<m?��F�7��t��I0���kLdr�~U)`s�E� Ѩ�{���jIɉ=edXʓ��.��jq�����Ͽ���xH4�ڨ�1��p�V7FO%\�!�E�̑�1r�3`4/h2��������Um��)�R���ߢM�_�}�S��Ҿ��kbN��[�T�>�-/z����ђ'j��x�Axη_��Ʋ��a�a���^V㔳f$�h`��׍�����q%��jT�L�J[d�t|���*�z6'�db�/(�'���d�d���7�`:q�e�R7޽[�ʲ����Ҧ'��N��#m5"9���0���ߠ�\��KzG���G�Q���F��b��Bun��Rq�J��s1'��3z�(8b2���R�`oX��q��
ὴ�k��Ϳ��?o�a��\�3ct�a��Ez�/�P�(4���5�S�7������]�>�V�T�+�Da*腡��̊=N(��&��8<H���Mdޅk)�n�l|{�������{~�����[���y�X>Y%�����Ԉܯ)�I�\'I<�Cwv♩��BN�����b�ĥ�]A��#Rb�6���[0��n^�
��r���@�)tnӛg?�H�{{��I��/ͺ�`T~�ۖ
\ڮ�-W�|r��,핿c�X�哗~!���nS���ܼ+ho6da^���4�#��n~O����K#���`4%��溧�8�Tm��A7փ*�5yFV
[����Y	i�ya>�ˏ�4]A�������Hp��i0�YE�{��,4�ڗHf����LÈ��;,�� �J}+OQn>�gh��xL��X=���{j�+#��ry�]gՎ�rO���f��BF�|Ԍ4��H�li�e���%�;7�cr*��疝I�W�or&�8A���+Ku$;��7�RO�ao��lr�!	�|�d5�몮]y�ѫ��d�C.���;N�'w��l&�v_��{�K��f�S���/����WI��X�r?!=dM���X�i�.�����I^�.Hg�X�9��rY�+�S��T��g��L�wc��EX�MRV:������lr,�.��M���3N��W��t���T劷�/߾Q`
"�%%��S�u|���{b+���/�dz�6ș����ʓ�
�e�T4�J60ٶ�$0F�#Ll�C�\��^a�,1�'tҖ���Reu��mn��mޟz�M��od�7)�klu�~��_�X��4/�������p�D��u\_z���I�W��DX��HWl��rto�o~e�)�lh�96�$?��F�^@����م8/;�ћ��\�k��r�<�m\f�y���'C�*5;�:��7I)����
qtY^�v�X���<�� 'B�1�V��w�{s�e+�x��+��TK֣�v�e��r,<=�$$$�#�C3W��m����^�����J��UD&}��������Ok񬎑����+�!�dU��Zbo3��������U�Ӡ.�@Tп���?��n�������?Y�n�w�i	��pI�q*uv�*��	�l
M.z�"U,l��c�l�}d���6	Q�#QHv6q��.��Y�daN/]%\�k�F���[��:�$�K�����Fn��Yh�b�F&���.�"޽,q��#DOm7�k)���6��Q+�L�(#��(�Hg\y��VE�H�S��'�?ޫ{Sȁ�I�S�F�n/N
��&�Cf�ɷr�]��a�_,U"�^��Z=��r>�<+z%xr�X�5�0&Ȳ�����p_`��.(��o���
���â?��2D������7�V�/�����_�ܸ)o3k�n0�>���W�8�qB�Ιd� ۆz
��	���[o�T�UK�o,��ׇ�v�������W�,eb���W
9X��%�b�aϞ^�"�(�!/}�c��&��M�7.��|n5�?�F-�E;�b\_�*�蚳�5.���p�=�2ȎR�ݝ������z� zk1-�y?�+�E��a}
EC�M�'�n�+^��3����h��hA��ُ���>6#[UR6�9J��D)�19�<&�kC�� ��ti~m�u
��X>�]:�mۏ*��_$6S�9��?���=�k��N�+~���o���*�53W�ޫ8v��L�P�с@,�����h��jج����
`dq��8:�s;�=D/$的<�*�����JTW�y�V�* �-��1�H��29��M��(@;���� ��4]���7��w;v�,	�9��}��p�*<���p���˛K���89�����u���7��I'_Zjn����ʖ��������$+{h����tBI|Lx�ى�r�W���˔�P��$?!]=���MY�F:泰�2�>� ��Du�M�tb�rr�VnKW��S���,ƕlUفD�GS�;۸�&���������5�5�h[H�^Q���O�fMO�-J-(J�ƽ��P@ (p����ξu�V��~5c��/�ˬ���f����v�*w�ᬩS��=���}���?Y�q	��U֗Wg45�P%�Z����]�p?�����Z�~	���i�y#����(�~�y��K��^ڮ,HB��H�9�|?滹���s~W=�m�$����i��Q�]^5z�c��V�'���r�p�^v�5�z������>��)��|��(o'�wR{�o��8��IИ��I�r���ξG����u��ۼ�4�l�0�+��	��eD��=@���V#8w_��?*��_���7��ųr��0�������>�Ye��WTo��x��1��%�� �(�`�z��/sI�D�o�V`U��3N��쌉�u���5���ŹĄ�?�BJ��~���ؕњ�;2��Ns<�Z�y�i���r�_�)r�~��n2�2�SC6�$җ�b�����t������(�ו��0(y�k����덶Z�H�
��'�K~(!��]��-�h�(�I|<�㓟��H�$���{y��j�����-CȄp���[���Ȃ��"�>����SX�\�����N*Q�ȴ����b���[؞�����]c;��I@O�����0�̭�K���Z��&rٍ|�JXc�L���-�<��t���L��������8Zۤ0�y�~��"�Ef�ۼ�xc��r��<�̬�ץ���q-�(��\nc���d��I͟z�4 �8C��篸tH��/�AP>�ii��0�I�SWEw�������j���(	M|��+���})Mr�\\�\q�}��ȝ���d:�{h�V�.�h�cx�#\��b#����|�+zCB�[+Ȼ�>���W�G�u�LT��)��_A��@�|es�n/�cut�:'|���Ǎɺ8�~@���zP�j��ρ����׼�O�b�R�c�����Y����	�o%<{�|&Mwo�B��|�g.d���(6 �9��i�!h;e��KbM�������"�ک>-?����t���Y-�=QQ�4����iN��7�(b P�s��ݺ�����fe٪��h����H��Q��ǎo5�6��^�&�)�� �e*��.���6��OҨ]���0��#b\� �1���*�?̂�1�oS��ϫ�?RB:�.�k��yR��[�s����=��7ys��rj�L<풐6u����zn�>)�SlQ���_�[:����uq����������_�,���eH�TB���.!|3~�������e�SB<h�`?��*X�7��3xD~;{�<�M��M�0�4����/ �qdޟ�ؕ��W:�'��ZIAϙ���hh�����2�"?n/�!#�������Ȅ���>�ގ =�- X�է#u��_EJ���c^�r��wA�	�$ê�>��J2�.)��L������`����l8].�֪��[���7��W�����k!1��v�u���X�=�{_'�X�뷓-C��N����g��
�U6?!�Z��3x�&)��^'�����xFv :�/E]��_k�\�������S��>�9aF`2�Q&i���_�-�o��mR1KS�5Сٝ�	�|����lO����r��Xu���>j;}�����G���tBE��	�hzP�7�@�i����]I�]K��F��̭9�W7��]��3h����}��mKww����SE���Q�w�/ۉqv�\K�b8��è�52��=� �|������Ƹn�w/���hD���	��x	}w$��MG�vko�Ę2m��7L�t���ӿ�Lս;�t�RK�&Å�t	�I_�ʹ�V�i
��������V��x�x�jR�f!��~��C���̇�q��0'�������a+ϳ��})p/���U@
ܽ���<�
b{ �V��-ZB'Y!�w8�v���A"�p�T� �D�w5�+D��g�[��۽�Phཅ`u�Ut���T�'ٯ���- $�K�7)���8B?HĦTﺎ+�
����7��Ueܭ�?$���p���~��r[�W7+m����`�ω���@��4��;�ܚ��8�1�ʅ"��v��^.�/1YAA:�6��|:���

�~������Ns�S��gϺ#`"%�/�� E��r"�v&^��?~�c�_8��,�J�>%��.�q�����Ϝ��]�� Y�-7��^���Zz.WZzl	��ȱ�\�b��è�uC���s&�6�� ��=|�R������@���
r0�lu��IF�?=fb�R�� � WzH��JV:7�E��q�W�&�Rv"v;��;�3����Y^��<�.��(��@�䂇�F]�J����f�?@w��(N���k��2r�_�� +��,�С.�q~о~���V���fN�6�����NG�'ci����VR-`㸫���te�Wg"upɣ��Ke7�ؽ�q"W�,p����ʽ����b}�k�H� ��C����\�����wo�Qf+4��"�-���K;5��tq���c�J�|�l�Q���Y����t*I-H���zO�l+K��h�UB�c���ճg���\<�r�rS��}�H��n	n�U��~����b.g.��je�B�F2b�?��%�n�\�tV��UZ�@tP�Rr�ټ�!1 !b&r���Aů�>;�ܘO=�'�_<��p1�������ݐ!;ܪ�vn��80h�q�m7�����>��!lW��kUk�<̣�b,/v���`��S[�:G+��P���F'w��c <Z.X�f6�`1!wْ��Td�;��O۠}Wp�EC�~U��ݲ��UE��z��7��/�?M�M��El���C����e�� �� �|8��!f\��ʇ�J��aѷ+?����M� ���1U��EXCsপ�����;�e�Q&)}��m>�w>2�q�����C_�P-�5Ir�]�o�I��[�!���!y�ڵ=_iқÛ��w�Ol�VI\��[���&��C]Z�;��=������^С,�à*A��>`�?
����Ʈֱo��^�+�.D]L��ȔM��C�*@���G+�즶�ǒ_�.�O��{}���u)������Y{��(j�c?���u���c�����S1���^���W�ٞC�ղJ"^�6����[�����J�2��z)}`�j�y`a��4!�ck�6�b�]�x�"+{-A��zNr�"�\`2�}u����Z���t�\��k����i������2\����֏.��	�����r���������|��}�b��8xl}��u�
YNԪ��_B7�(<�-��;�^Oc��^�������O!��<uD�C������8��hB�``�R?�Ҭ(@���q�}MHh}�W�δ/띜o�u�U�+I#�� ��>rR#'��#G?q��<G���Kt�ޖգ��8U�����&��^.�C7����H�PT�*����7m�M��X�a��x{�����w��o�IFHl��t;���qd�]
C>-Rg�.ebe;��D�o+N-/OE�m����m�Ȃg''�3��v,��0Q�U%��6���c(lb)�5�ϬXBF	�.Wk��C�!���*A�j��č|P�]=-���^+:�NK�T�#�]�'���q{�d�L� ���VN �����>=��*pc���Dw�o��	��0o#�X��<j��(�A��B����U$0C9F'���ǝ���u�jO�N/���rYyNɑ-\����Z�d
;��V�6^דv������=!�ǝUȔRW._{��t�C�ֵ�/�z����#������Z���{�.���<M��*|��K|Z�ՊƝzI�B�<k`I`���wU�7Cu#3�%P~��@�XZ8"�M&��f:v���7�Τ�;m�������!�u������]2G�I�g���+���E�+j��t$��{*���=ۮ^����@ł`��Y��,�s�@���}�B�� .���������v�nB��5X��Ωg�9��*Gi�{�9fd�zt0[��x�`���ê������ȫ[�X����-�Rv$�Θ
�����_�H0� Y�r�_���X�D��ݻ�Ϟ���(k��Ctө��.�)V��3q�uEʢ�f��y����K�+>����]���SQaR��KQ�t�ʇˍfe)�T}u�]�r���`l�ٕ�����Ӿ��^��ʗ~���㮝a���c��z�xX�,_n�[���ss������A*]���8�x�m����7V�ը���?].�3GBbJ&'��
�MQo�Hh���8�}-�b�n�O3�ʙ
�4�>�G�̀m��g
�.��H�):=)5�c�$L�����j�tS�f�R!P���#w9U��zNlU�V��&�ʖ�/ŧN49�����E��+��;R���nE9f�����H������:�"�5�1M�x��Ѣ�6N�Pf��ߚ0�V\����p;���"ʀz���m�1����_���Y�MY-��{d�H���x2�v�n�m�4�X��s�������-W��n���9e��|�������.T�k�;�O,�[������o��k��z:�?{�m��YXR���<��K�x]�e��eɛ��s��r�u,:̮��)�'#�E��^��J�aųgTd �`�^ǻ���Z����D�y�`��sz�ۣ���g���`�V�"��Gz��ꍼ��̃
a�!����AV�Do�-�j���RPǱ��}���5ŴiJ8X�5t
E��&��t����]�R J&��eka���.���.e,r��X�2RօҴ� �E1)%�+*{�����:��0F��%r2��-	з9�7`��A���6^���f�-��p�$x���:�*�w>Yb��b��"�4J!��30{���L$GTF7\�e�JE��z}g�A,�O��L�f&Vd��s7���/����c�Ў�Ȇ0R���:�2P�y�����7�Z�&�j����
��������i��S�`_%I
xRC����hb�l����~^~N(!�\�|��ߡ1��×��A�^H�>
Q�?
�5ղ�Y����/ 3|�8�
MQj
�?�wS1Ў6��Nme�G�҅]=+�r�.}�d�CE�bQ��������0���/��S�o�񥚡�1R����?cP\"��79Tc���b)�M�k���ٳ#g`�q5�8D{�(��S���Gps(kDF��]U��C6�9�+�&+�ψ�s�k��c��0G`r�U�=D�ִD�^�n'��-\"��?5��>\��0_��N���U�ږ�ls���E��+�K�~/��Ŗ.��O!Ҟ؎snc��K/�]� ώ쿾L ��p>�Y7]�����#�q�f��O��	Ӓ�hJz�e� fW`��*�� ��,����ʟ�D_
^# ����Q�_�m�/�v]�����X�82�Q��~�f�2W�'��^@����������ޜ{u`�:.��i�z6��L��
�w�,��U��!*'��%,����]�\�{>ԋ|w�}�Bޟ�=���9. �ݝ�-Slo�+�3�^V�9B,x���x����d���5z_-K{��lt�	#J#O�ٗ�����e�~4��v9�,B�:k�IW�6����r��k�voل�*A[B^�b��R��v��e�o.����N�QV�B�,T��LF�+��u7S�QU�BnS��ߏ���nɅ4{۔
�=Tƭ+�~u*')�W���ͻ�?�m׉kb��`���+j�yŬ=���r�[���3,/y�+q����F=���T��J���3#!v��(K�m $��If�8���L�E�([J����[+S�����
��8f��޾|��-���_����a�ź�({:�(q��D��h7?)��ЬtR�9��V/�%vcZ8p���Jf�r�O�D��q���m���3���)��;�_��P�U�`鵰�u��n��l�����7�����zUTR�%�?kB&#�gݷ� $;����xX+W�ʗ�AO��//���Xߕ���p���'A��]M�	���~���q���z+���{#^��h�ī�g�����Ɂ;͗�%�� �"*�.S.kXki���Z�1��*w���-ъ鬌��P7��"�U�,p;����h�<-%
j�].4h�<�Qh��- ��SN�T0��Ȥ2csOӴ��V��_�E�z��6S�SH%�>�&�� ^h�ѻOx���ֹ�|�&O����M�`���Ų�Y���߯�w��C�}�be�w�yz�E��"atP!`L��P���Oυ=���~������c���@���R���o�Y	������r���X#�6w/n���D��pL�v��f�8n��I+�fh���9�㉦�鋯�x3we�/���~��\kR�@�<��$�|���g_�+h�ˢֆ���9�g�?�IXQ�R��������1�%������!*�t��_޴�L��}�(�l��'%X���;sBx#�ޝ�^豬�'3��T��/(\���P�K~T-��Y���y������[�X�
��]��߸إk�g�V%�����S��^1X%��W�}��<��M�"B�p�1�s���i�x�h���O0}�c1��{���b���@��Ǳ���6���E\`0d�\)mqF��#�f�������4�����ZǲИX {j��p�@���ecY*덾\�}��<�T����g���[����9aa�y\J��U���(�v�W/k�,lx0�.?�%��|Ų���gMZq����e���0�$$��2e�8"�;"�,+�-�P
������a}{��C8%nr?Z���� JKN�S}h���p0S�������������{�)B�^����HEр�ۗ*f��u_�V}@��x識	�� E3n(����Y|����nj��!l�Q1/Z�z�4~+�|l���4˓��n�qKe�(� �Vd��;��S_���iM�"���v{��=ܬx�:b�g���by�I.�X�n"_��Y��)��?�`�Ih8ǼN�?�#l��i+]�,�,�~�9=���)���b�w����N�?��K�����M��uO�L+�߇���Q�g�:)�(؏�+�>��/1m#)J�t-����iTe�˜:�eӉ����/��Aƹ5��ùF��}�Ug7Q3�z�+ݿ�}1�8�<O^��C[�w�je9��A�y<Z#I�Wr<pTe��B���i҂�ʵ�"�UӖjyZ9���yZʄ������gh1{��{aO��R<ER�c�۶�~�:�����2`+�}����]��HG�Y���ݩu���}Y}&IO��*+{�޸�UbX��x6D�V�ez��"�-�$U��u�0l���l�̛u8���)r�Zس��"j�E� �a�O-����q>�T9�w�>?��@����LL�q���%2��n?��E�FF�a�͋�[�VE@����O�'w0X��KP�0���I�1ο���G����z�I_aծ�����"��2V���g	<K�#þ���޻�|<�ỏ��}�"FV*|�]WT�V�����t=�d+A�O�i�:���$�rƪ��H�=8��h
�����teV�j��pE��fz\�Խ�n��3/0�w�J"��غW4��~�B�eӊ���f"
�����V��p��Ɛ���H�B�#�P��[��>7�����t��x��m;��ن2�ޖ� u/��KBp�)P��,��B{A��5��醑�~��ݛ�oͤ2~$�˸����W2����-��9�cRGö�����@�Zy�~����������'�Ӧd6_#3��ϗ�^o��	Y��=o[�ެ��q�;b��tQ�_��Ɖ}�+��DP���U��	���^M��PСZ2<�k[)��؅'�Y�G�1m�	�y��q*�_zu�=E�N���o���A_\P�1��3e)���=��N�^�.��r>(){~w����`k���ȮJ�YxJjWR�i.���I�f���f��'��VwYs�:ShT]c�;?W��g������������x���`����O��U"v>��`��wr�S�&r �L(��T��f)�o�}��޻5s��/,X|�Yi�(x3�+�JFfωA��S"�}�;r%�g�?]�Hq�Al�hĤ����tjv�q|�P�{�g7/�Ko�,�<e-t{��{$�y��5�����틳�%�YԎ����=mc�ޢ8�#I&�"��?K5�E}dB7<W��C�*����Z�8[��v�3nV�B,���&�Ϥ^�s���ik��*�H��ў���L���+��|#�e`��k$}�}�Ӭ��ìŶ�$J�?r�}iɅ�*��5���������3���_ƈN�\J�]�f�ef�V�P˭��G��`nE�~%DmQ��P8r����ݿO�����$=Z�o�N�MҢ�Q��s�
��^��V��3�_��~NIs�1*�zj>��jى7�W7!�ui�ݘm(�|2����� B�i�[��s��m=����t:F�߫B��⛤��c��L��T3T�ϫ����R�v)m���?���� Ga��f��H׾��ʭ�)��rk�)J�^o�f��:�F�n�	�H���Ӗ�����ػ�Z6�,la_b�D!��ɑ�5Ы��4o��jHGL�*O�0�����S]������>�~��J��+��"��w�Bg���WS-R�Q�0;gY
�P�O�ܻ�Iyz�ZD�z�aQ�����2k֮(��H�=$������Y��p��@�*���/�ػ�v����"{ƾlj�P0������x0iD� ��e*JW�� ���*eZ������ �v��74�ʟ�Q����N��F��g��p���9�<�ߤ��a�ؙ��Q�!���d������C��CC�$ۼ<cb��V%w��y��yK����u��)�Fuǅ ��O�N�n鿅�r��J$��y�Rՙ/���w$]�	���T�%���Q�߂3�+��s����Sz7]���0ePJ��7ir�0a^�Z�{�!�tE`N�5�+���z�@}�I
����5Ǐ�RW�������V7M�����=�Nh-�dİ�_�(N�Z�E}%|L;�
�h��g
�u�GDV��y@�P�v"�7O��9�~0Q�J���N�h�ӴM�B�8��ۖKU2l�~�n?����\xդ"@h
ކ+D����Xh����[.�=��W�7���r��|#��ja
���6������Y=,��4���;i�?�<�w�\��"Mr�s9�Si,"���v��{�M��Il�\o�S�!�N@z��� �V#���/����qj�d�B7�=n�+���극@7t���������;9	���$���(���M���a%�ۨ��Fs�5}���b��4p@8�5 �����귫І���_b�ث}Pm1���]	�0)︪H��׆��?i�D#�Ǘ�
Q��Y0h<�y��Y�)�SQ^` �����-�Gz��pʺ~�$��6Sw�l���1$ +��zE�eN��b�5��mjA3��f[BL�Kw�F7�*jU ����[ډ0U�-�"0�n�B'�ƣf���=�N	́�Y����D�I1�������:������nN��IZl��N
�?�>��Td)� ��/�*;�"��ͫciA��SlՀ����ی��U�*����*MdM�h�� ����7jh��]S���=�ws��+,�3���/�H�N���&��p��p���ti���
��¿|8���f���@�0���>N�
��O��JC�����8�G#fT~��*�	�C�4?�� m�A;�[�)�_F0n�h�!AT�m^��` �t���r'c��I-��2���?~W�jOi��l+ G���J�ݙ�la�m����p�Aİ��j14{�����,͒`�5�~n"���_��i�����1�,J
��6kp��k�_a|O��S7(�N��h�	��BW�������3�z�L;���q�hq1��)�Т��@ZQ�����Y��0��W��ldG�D�A|��5G�]F6Z�?�f�o��t��2c��>U5��>����_��9�-���%)i+�X�OG�O�Z�P��D'��T"��g�����TxM�b8���٨�*��F�<y�hl�.�-�#�9�J����w���_E|III�}�ity���2��T"rJJe---�����/>8��dvS��"-�(�1�iVI����k54��uQ���)Z�s�5���
�;����l��O�����B�0�.�
�z"�0<�Dl�p������y��F�]�wп�����x�Ȓ�4��d��5��q����P��8���`���0�b\Rol���=?+a���X҅ �u(�F?���8�����_
��bV��j���C�9�]E��{j�8�r�q8���GԴ�������W��;���2f:����;��h��ќ����;UQ��<^�����y���4V��#w�!ײ��2��8�,�����G�T۸;)[���	��ꨈ��ƶG�?*"B�2����֢'�Ջ��v�a����Ш3�Z��|�*��������x���S�V���&Ԋɢ�K�����+��F�bX
1�cc:~P�Ѥ�o_�l�v�&d_����^��^��E��PWJ���+�C��Ȑ�!���1����ii����)��B����Y��ֶ����_d0��B�F�0)֘�J�_�5�9�)�
������`p��7�t.��{{U.\ �p�f����H��U�(��G�����*��D)]Y�sz�B��6��[�w~>��ŋ��W�����yP�1��P����+��i�9�Jî���n�8��{.4E��P�ɷ-��>x\`o��j��~��=�N�� B>&8��"@�J~���_�=�I�2-_nn���V�R��Q�`|�x3�eg{�o�"g`p�3��,O�cU�qS��a&�(��P�D^����^��~�ҫ3�L�0���ٙjM�����R��^�I�|��blwW^���������/�x+�\>�z[̵��!��i;���C��Z�B�$��ح>'ҕ2�Mb�k�c�ga��ԙO���5����+X��D�m��}�h��`�Ì�f�M8[a[娠8/
��)�@���q��&��L(��q��(����maj�/=g��V�����Ԣ�s��^���Ȍ��S����_#"Z��#�AĮ� ������?�~}-+h�ͬ��{Tm��,�8[-$$�z��o����в�c�A��!׸}�5fuC�T���O����m��33<��LN�N�s��=��1�� ��#�������p�Y�߳��1�@u��?�d�N���ER�d�睡��s����E�]ǽ7;��ݼ"�/84�����Ν���Ȁ��L.�ɋ�Q��n14Q�v􉍻���ލ+�i�����FY�y�7������w�{�'��ee�g"Us�֚�����[��B�Y_��K���-�p}��]���JIg]��%<��o̊R;gM���4�^*]��s��i���]����W7�p������h�a��j��=s	Q�шg��ޫ�9T�,��b���8}�[T/��$i|T���VIi	��k|w���Z#�M�&Y*���boo$6J:���;7??2""��˩fܑ?I�a:F!;����ffV�+�L��J`}v���]~���!T��]9�T�	ɢRfFƋ���222&\��Ŵe66>�׫�l�lni�`+G�^��f��i�fuS��cbf��eP�(���������ˡq���9�ȱ�Rq˗�H1��o>�����;+��(�x��"�˃[�𸘘�����TTQ����9�rv�k����=7~1nw��2-�t�f�Д����V9����{e�{ص����h�U�2���bhi�i�X�SpgmQ�m�^AᶒV�%+����ohߡ�@��h���z-�3����O�4%'|�'�{c	�$�!��%��-��.��jVP2]y�o���z���@|Lɻ��X�{ff&q3�*�'�J��X���)�U،"�R�Z����������!��T���d�9r� ���7�����(�H�(UQ���g����v]�qq9�B�����eB�-��y���Ř�_r�/�<9�Ⱦf���z�5�����l����/ �ٳ`��@N�q�q���y�{{.y��9 ߽,����Y�V&�_!:�C���x���t%�Ɔ�L�O��fr��ӭQ;�=�noo��`_�{�����$~�+��"(��5�����W�%�����kS�D����۸a�U@E7�����Ł�+;8S{-{t�Q�Q��ji�|)����P4>�i�?��#�z\� ���d���gfeU��K���,��Cxt���~�vj��IQ�kjh�KAЛ���a�gw�b�V��A�
X0��
S�A�sǰz˃ѡcZ��c
�wl*
�E,rd?T�M�Ё()y���1Y�'W��o�f�T��9�����働t^bb�
/�����
����ڕ��^-� R�4����"$��v,@������x���Y�������Ƈ���Kf��K訠?�`�qe2a(����uQ��4-���W��~��������Cu�o�4*6����,���"��J����-<��Ty�p�r�+墬������BL�/W�*�K1
���=�<�?2�#ޫ�l+Y��t���>{D�/6��%ך
��zV�(?�t��#e�!�B�u�L�5h!�3$�l[�{h]� sM�$el#w��m������4Z���Z����T�0} Y�.��qk������ }��	~P�L1�<AI�uwafc����J?8�P!�=tH�Z'��MC���TUY��>�J����\�2Īƨ��D�	h�_�E~H�
z��ݯ_��dq7T�Օg�>�^@B�룅����?P�ػ�� �����K�?��&��0pY��a@u���,����{�/��Z/�B��>L�mֵ��v�]�.����984����V�B4#�m6�i*�ÔO�p���%�����(Z��$%巶���E��v\������%};I������Dj&}^ ෶X'��+W���vě�<��(����S���L��~��{��1�ˮ�e��W<����dA�*��vrDC�
7|~�� �%�ٽg�_��޷wM�?���/]}u\T]-"�tw�4�H
�)CI*�]"JI�P"%  ��"�tww��w��}����7p�9{?�zֳ�>w��z�u�?g�h�mk~���d�H"Gr�T�?S�YPk�uZ���&����X#Z�av�ve���"����Xw��d�^�:�uu�t��k>̄��
�U��%g�����v_
����]p !f��ى����2��_�?���\��|x.�S�(4=]�C���=���>�%<�
�U(��G?:݁)m*7������vz����|��Eod����2�iXe�#��Zq{ϸ*ٽHHmS�J���N-p�����ЌmM��w:�<��xRE<�|N��j�/�%������U`��*��C(mPߑ_�=���nҶ�����Z�_�!ۄ�/}�"�S	D1	���0��-�B�l�}�at��;�5�J���T�2����QfK�w�C�r��?��}p��g�%�:n��o���h>}���ͽ�X2�Ϛ�j--Mz���f���7�~���r��=��I�583	�Δy�Ejzmgn��Ћ,����|<���Ζp܁��Щ������R�|O��n�f��&�N��n΄k�l�aj�'6h��A��4>"�J�%"#���S�A,r�7��/鴺-y\�''�w�oT��~��E���޾ɼ<�_�?W���!*����/O��%C97y��7|���K����k�~L�҅(e�8m��i���M����r��-�[Ai�$6��k�?]W+M��L���8�/�så=��n}����,u����|��W����E����p�W�i��??Q�/�T6#(��h�ْ�R�JG�;-�����5\�e��ؚHJ���}�7�>V8��!)NlDa�9���3C:�ή�>�/�� � r�@���$�&l�G�ՙTooo�p�ZoW�:C�m��i{�HL�k iw��^b�1o�c�Z
�?��x���92��=U���x����c���P�l�V�tdA��ȝ�$��r�{Mjx����6IQ9�WuurR��~��>������}�S
��`t���!�Hp���A���X��6a���d��H�7�Y�
���$b��y+�����j��D���)��+YLo�Y)!��g����D2w����Q�BF[����/V������t���VO�f��#"���}����8A�T��g�U����#.m�郱�>��@���57��j���Wlͭ�.�6��k�j��ք���o�b�P�Dغi��_�����뀋��J�`�
��*4�N��ъ�:`;o.3R��{�6�Fe���lw�Σ=)�H��1q�yW,���
[�X蠺�+����N���xW�b*��y���h��z�pi����ﺝ�AI�ǳͳԴB'����Mn���n��fx�2U��F�d��I_���Zhq�����*:�#Q4���.パ1�ݭѐ�LQ��)ܜJ���]_�5T��@ 4e�ld	�{���@�?�}I�ؘ��G8ˀ��R������_�� ©���f����h�4�ݓm�����rt���>F�)g�^ (A�BSx �Z��1'��?���ĲM�f��<��VDP�����9��G���?�%)k��r�{�g�(�x�ZS�pKĂ��sC���_�X`�C���ۜ_8��P{���mx�Z&�"�{_�O��5TM����\�`�
�8z^�W��x�0�����l+vrr������b<5�It۪������.��;�}��Z��v�o�\�e���Y[�~+��AXDt~|��fBt�8P�D�6ik�8��<�v�K Vq��T�^�9�z�V��|L��{���d�g�'̿�KtYQ�l��J*�a���ޮ� a��8E�^�B��3 @�� �	�����;L���G��c������gi(���MX�������AT�56�F?qX�z���A��<��%`�3B-y�ż�Q������j��:L���擇:��9�~��z�}�h�ZU���eL=U�{���.��Ff�f��gv���9�6��e:���foD\����CB��f|�N���*���=(O�!�~�>e�c��xQgsp�-Qٓ+,��ǳ|(&�OQR�O��G�ύ���r�q���9)))�' �ń������Y�=��'�:�APf�MBm�P:f���dS*>���6��嶯#��{&��l�L��D�啕� %�+���>�m�:��� ����Ὁ�Y���2s��������VM��Bv�;��Х��"%eeK�7��BAGB�5�	�f..�����L�Ԓ�Nu��u�^�4��gW�������������P̜޲!��Tz�}�ob��+��u�,��9�����:�}dF���g0aL�i��%֬X�ٟ�o�<Bղ��
�����I@F�y^fK�H�, )�V��Pqھ��a�V����-q�Q3�W�m��r)��%=�����#7\K +��94-� !�Jfhm��V4K�����4����'<��C:�m
���B4�J��X]��IJ��/U牚;�kc�d �̒r��X���Ub��̍�i�e�����*�'������F7L��&!��+.�p�yi�= ;$uSY�y�G�*=;j�b���$����2�(�́(�ql�)�����z����L@ 1�ݛ���)G_�����`��~2,�~�S��r��������mB�e�fl�|���Y��MW������fNŌ�2����V��sC��Ĝ��~\1bI�y���C��\��)�"Z%b�F��;oWc�g��#���t*�,�͕D:�H����G�yĮD��W�A�`&ϨO�z��#S�#�������\����W�� �lw����us�_�g����H��i23���9�П���!F�V޿�^��Ʈ����{/�Im��{ҹ�Cs��a�Gv��mZl�7�c5��3Ep�ZdogA��m!����ek�#*B��6|V����Nc��;�ĝ:A�+Zs�Y��p�Ą��	�<`��bdddM[e����m�>��94��T�U�z1��������_�G��x>{~Hʥ��WJ}�;`@iy����~���Ӣ�d����w~����o��X���,p�X���z�IAX���p�痣�?|/ҁq���d��������(��TL�[Ș�`i�6��u��ׇ�V���pݸR�4,��&���a�H!n��ͧp;
�>��2�*��׌

�4�Y�fJ֜�C#_v��Ơ��T�� Q!щm���î�m�*�U��J�-Xs+X��W��ٔ�=�T�4d�Gވ�k�P�Dޒ����(�Gv�=$*Q��tnr?��y�L���dɭ��v��]���k��s��x���׌��l��\C�^�	B��!��d`KPP�N� tXNe�[��M��������}�S�>�|1R�dlt4��w�ߗ�I�ϩp~*{o���Q:�<}|ȳn ��g!c�U}3ө¦&����P;f�ϳ�Hv��6�����A�`�2�3s����^FO�l��}E �6L�~傇������K�~�Sz���1M9$���8� y4��k��Bww���o���ȉ���?�U �[��t��G���e]�2#p�x����S�m<!�	��� �4��'tE�����kmV��;��Q�u`ya3ܝǵY����^�ٱg�lOT��/h/|�<�%��%x1�EQ��N�"a���YU�k͟lt���<��y�`+�c�ː��T�k�����|���USe������	]z�$>4�hfI���"	�W;�"�_����	��Q�j�cD5��������CQ����:b[�r6��r��M�1pw�!���l�a�����[����<�i�� ?V���������[(b8��f]�^�w-���&���Z����3|u��]�WT�����ʈf"%�W9�.t�\i��Ũ��y����oN֗��n�~X_���|ck�������h	�KZ�ռ�n��166P���r�+e9HZ�������:���ubf��?}�MO��3�z#��ж�	%����������
Њ�����e��?��5�O���6��|����#��Xr��EMC���W�7P��5���{"BCS����?)qʮ�$����Z\��@M�@-�����{vE3��gf�gϚ��/��pj*m��\o��K��e�D��i�'�����v��_(;�Ó�׏� ���-T��wQ������>  ]��8���2��nK���Z#Q }�(r��%��rJ��)��|�V�}��	��ѥ��ez;�mS����ώ��w{_�)�7n"����2���j5�sIh��ɯ�|�P�ܕvv�+Y��	���^�����a��Ә�ز<���g�x��SP���́�w4���c��sIa�ج�� -~��*�c�G�Â�Bo����{\&l�ؖ�੝�������V�����]͈�����'n��D��	�ͱ_�""��`���D,�1yr���*>Ni��l�Bڎ�D!�T��05��5�k5/,�Q,����6��D�S@����Q�K\n�p7wq�?dkFpD��ar��4Bd.�P	u������HL��<�T_߀�y&�͑4.�˟�-���ߙ<7ܖL`�滢���Ox��J?xV�HH ;п)è`��{���w��4�+Ft�4(D]����V�wVj��*  ����Ն�'��a-��yԛ�[�#a;;;��� mW	/'��:�� �Ŝk�j(�����d1=:�d�ܷ�[�03$�f�j&��C���3���8^�ޞ�8��ެ���`v\�UM���卽ۓ���pD�~l��g�su瀞4P_W��::fJ(-'�E�F�A�]�/�)����=�������ӝ)<�77�5���iH"u�?�4/8�SΝcd^��� ��uA�q�|s<պ�-��j]dx��ٳ��Uk|���5��d��mҰ�����>0�
�P(l���eb��٬�2���`>a�Ƃ�6qp��R�|T�VHt9���?\gMg���g@�kS�}��|p�G*N.uX�I�H�����Bwq���Kt�a��s^*��*�2
q�Iq)��j���N�$�켼�u�����j��ݽ���=�e����?�~�\b����iļ_%Y���{�y����=A�@dd�s������޴cM�c�h/��H}}}�ggc�������]�����r}����?ha�ꝡq���] ^��a��ެ������5P�ΰC�`�'�@U	t��X�7D��D�Z���~��.fNT"<ѓ�!�@�s���UW}��[9g)�uǺ�r22�����C��C=�zEv��ʽѥN�f���2j��L�� ��o}��g&wu��ֲ�Jo�d�=<�<	e�|)v��ZD�yD{�9"m�
#+��\�r�ϸ�w�
Et����1S6ZT���ڣ����͓�4��DG�R�z*�	D�m�=S�p�%�L3�~��Z�9���)n�< �*�[�T�)�[!����l�ht�>�H����rd�y�&���>A�ޒ�X$@�@%w�zAK�%�h�a���������s4�ڜnh}y	i���/����G��^�]��X��/����2�KV}��8-���Y�RlkYsӪ;2��<����L���Mq�ڿ?������|��t=yX�ˣ�L�7��]&۬�5�Y��5Ȗ����ܸc�ͤ�.����2%$�P�Vi�)f!m�ޚ��~M3�{�1-��ά5�#�]r^#��������D��`�J�X�y�N���A���آVc���qR��8
��c:�Z�P��i������H�9P���>�w�U�Z��_~�}�ts��\DWRj��n�����^2�2���*����4g;��GUp�zw�ߙ1m��}=��ĸx \z=Ǣ������c{ȟާJ�׆���E�*��@C�	����$P/��Bk٤��nkL�4�x��z��q��_������GP< DJ���i#n�i�
����k9���襳?�6�y �"��ōԦ����YN�h%��#�������0�^�_BS�\k�m�6im�("CaҠaa+�,"��	�2�T�,�BS�0�kg�c�
W\$蓙0-��?���;Wnޛ�9}�i��3�'r��uQw����"�\��d4���(�t�D�X݀� ���$9Z,@��&a�0��Hqcr�wE��1@����\�����%j�%b�S���`��%S$-�
���nc��F�}�ހ�ڢ�7h�H'���TY 0�I��N��0ǩ�yq���Ah^��R�5��*�^�:W�IN4,T���!1��}��Lz������E
��
C�R�L��@a������3�³��Z���b[�sO �(i����Bomd���C����9�9e��C��8�k!�W�]̶���K����H����)���ې��BxcU��l���Z\E����
���Mx
s��<b�(�'Q���:�O�c�S�_vH�3;�Q�jA.م�czc>�ﺳx�G�S��V�eAM;eSkQճ���N�"�0U��6ʬ����t�RGE���n�@���8���d�k�eZ"3�����ŝ�{Pf�z#7*��T]�Rf5���
�N�Yd�TzuX��
V�y8�F�.��w�dК��{dkHttt�����j���݀�b�'XX�s1�d�����0��54�It���TהԪ�	��f���g���S�R�ܣ�,�i��+i\����I���ճt�EPÅ?u'���*���ʖ����u�v��ߺL�i�Ԅ�O��ќr��gN�ecv�*�
n$���xR�Y�dr�>�_�"���d�\WMT�J,���i��|��K�·h�Y�c�w��z�	-�z��wM����ch� �k=�g��~"/V$�=��/N;P�E��|�R��tG,�N�@U�X��u{#_��E%�5:sQ���6+].��cU�
vA� �a7>fm���n��~�B����]ה.�!�y��w��w"fMC@��Z|��M�1��޲)�T�����H�1���Oi�g����r*�6��'�O�M�Jw]&�~,��˿h�zΥ�mE�Cz"�B$��������Mn�"��?Mi�â=c�J�fҬ_�n*�p���� `|�jNX��Gv{�摙$q-w����h�[����f��2\L�q�]!%��r1�:�U%� 밧����ˤ(͜P�������w
��s�dz��zf���O�����4VKq3�b-V�N��hߣ,�B�UH,��6i�>`��ט�sL�z!V�RgW���m,M,c
U2|-E�����	�1U�$!U�sŗ�tr�KwK�+�6�Ϸ���ې�cdF'�G��O[$MwiOȫ̬ʴLC�ph���t{"W�""BAy?��^����E/샳%�B�6��=<�	N�=O-�CtJcȉI�+P�n{�{�V��^SI��.��֍3��m�U+"���,5�	N�98o;ɯ,������#��U]��k�h:�2�Vr���^�uO����*�T�R��ˏ_��M� ����\Dzo��E�U�p7jѢ�D�Y�B�g����^��D�J��fO�u����]{"�a�ܴB�~H���MH��jI��뤣آN��4Us�b�f��`��9?4������W��m��4ʇz"�2�����bi�
U5t�9>_��*�b�&h�W��nzR.�:�4D���?F�!�ԛ�V��yo��ĵ/1��$}B����<o�}|�m��:�
�t�Ħ�mJ���b*��O�|��Ut,n�#�?Y���	�L�ɯG&�9�YM~��6�cv�@�B�����z���� ��f�c{��m��Ͷ��170�j�}�OD��O��o\�MplmS�.�勬�o���P6��'{yox�{������(��Z�.�u�z�s?Qd��TW[�N�������p�Bp�q�W��Tv�H/�m�����D22�9ѵ����&Q�X�mBoFs�X��*J ��^I�23ۀ���P��8�z%&��@�\�o���]�_� x�&��G���i�����J6*�w!���1���ә>R�޼mbK��:m�]>�Ҍ^4��:_#	��tC.�����P�db%�*��5���ǥ�`%��B�7�����c�ۯ�̭_?Q�]ŗR� ]���xP����B�߫z"�ˬ"mL����~T�MwII\����9�n^���?F��� ��ݙ�o1�VN�V�6>�B��m��������&�3'5��k�i�왕���4)vmH�
3)���Z�5�g�F�2���+)�+�Ӊ|�3�o8e�Z-�3p���s6J�#&�z�ٖ�B>f�֏�u��gI>fI�SS� ��u&�(�N���s��M��|{�	��HW��_����a�<��0�>w)F)�g��B5�xw|�&�������M�rV:�~O�iv̜�N�;��I	�(E��bTp��p_=��z�iJ���]lؑ��޳�V7�k�����{��#��� '�mJ���F��`�`1؃ׇ7ח���R:��;v�Z�Ab4k�=��6�3�w�~"�L���/�y�f67���ÂB�+&9���{S9�B��{]+3bq��1B�xC�ߏ�cx�˺�ٺ���X
t�
�ܺ��uJJ��L���QyQ�mr.W�*\9��}2��(2�n�w��ݙ
��vcG�_7ڑʿ���D��̢X�U�+I�����_��S�|9�Nd�3J���
~����Z����� a*�$����[(�����$],�~:ř��~|rِ@��O�%Il%�����C�EJ&��B���NBx�)�VS]�DKi~��c(m~�� �Ĉ�9q+'b�$'��ن�-`�	�����d����yS�ǚ�S@�ʽ��c=}S,PB(�5&�^]��1v�_u&���dd�I�i���Ӻ·$!�d�.�q�.�j.���,ۨ�d�U��C�Q��?�q3�Zo`r�0��/�����|��)M��t\��B�c$�.Q.ͦ�d�6i�z|r��<��-څ�-j�~�fe�VUxs�S{B]c�����������\�G��#�1���3�����H#���7F+�=�Lʲ�jl��/�572��\�.7�N������!�ZD[[�?Jw%�'_�!��)0)���>Sb�䎒bJ�����)O&�I�
��c�WrG���,�i^Jh1C�I(�bQ7!�|�F��Z�*h��5��n�����}���w
6K�����s��i�@�'�߽�_�\����'�DQ��D�K�I�JD�xI�<�~4�F��=�7O֑��l{�B�PO;;vdD�,���5�%(v�HapL�M�8�Z��\�}������!����xy<M�R������a�������"*
	X�оNLN~B{��x%��Ww��7pt��(���8
��(`���	��y!7����{�O�~��ǋD��K���멽���$Sin���]��Ck͇�cJ�6� L���rA��c,т}Q�9;�����2�\��t�+���?1��e7/'�����fTr�1����tJ����iE���8�{f���v�]1���c�5��9�)��"\��GıL�'�m������]�M��d�w���{�nO�I�p���d>�������:r�f��1���քK�Nn�ԉ�)�UCib�����,�/��1�Bsw\뉬��%�$AX�V!���cʗa��| �Q�ѯ�!��/)���W|�����L��� ]��w�uO��yWz#�Ƚ����v��VF̊�N��� Z����G�y�X ����g�lX�&O�HR�:p:�ݻ@���O�R�e>rj��)��?���G������*��"��h7�>���R􊨷��/�~��d�UЯ��D��B�Vx�@�G�ٝ��
�@.��]���Lv�Dl��{,,�%������G�!�B�~+I�`���S�wg���uvٸ*������ڃ��9m�he�wL����O'�N��HT�A��8��죞�{�!t�������!k4n9?���,���Z3�À�_�}Ԝ��U��o�?�H�!��$���x��-m��A?�"�ݟ�+ʪɔJ���PK   �x�XQ//�@  �?  /   images/f7eed1a5-74ac-45f9-b2e1-80b6b3a4cd0f.png�?��PNG

   IHDR   d   �   �#    	pHYs  ��  ����{]   tEXtSoftware www.inkscape.org��<  ?�IDATx��}�dWu���+Wwuu�=9hf4I�, !��$!#��l��:���v������dda� $��F�8#M��Ω�r�ﹿ�����C�hhy�F��z��=��}��?�J�\y�#�zy�L�C^�m�~���f��y�e�pM�tY6^^^^��]�]p�>�&��Ws�o7�A���a� j<"��B�+��j�� 
p����&��qۃ��A�2��W�v�q��M��W^ߒW��
�|�m��z+��_�wNn�	@AD�7m�tg���Vc�����6=�`.O!W1ö��D��YOIo#�:�5b��/Z�x-�`у�t�
��8�9-�!y}_^% �a0�􅢌@�q���`Iw�E�2"!B�%�C*�	^�ٗ���Gqi~/�'��f��d�l�b��x�O@�O'%C>���:y�A�k�ۃk�GU�w��:<�Z��s�����-g��FM�Q,�j#���=Y��)t4�I���]�e�X���$��qي 6ԇP�3U=�Y���x�h;FeD�]���"+]��._�_xg�����a�qd8g(�ɗs���(�^���?&���=�+���ʰ�ӰW�����t��"��X0E9��KcM(�WxqZ���^�h��ݣy<џ��nӭ����V��lr�|f�yn5.誆Gv::�i����ޏw���\__y)��i/���n���� n�SO`ݡ�`�ɹ�H�]Y0+@yƽ8Z�r@��]��zd ��?��W����u�v<�n@Q!5f��΋F�Y1|�� ޾�U^�>v�KWظ)S�O&q۞,����wV�06xc��K�U��Duu5����)'1�:2���8.�x�*��_>ǋ�B5�
��ߋ�N?����D>:*h(�|}���Q��؟�=��?.h~�\���yؑ	��1�ʩ�ş_ވ�!n/BUU*'�۹�)�N�L$p�f7N�K�Ϧ1T��Ja��9կ1|��z�k�C]c3��$��`0���:&0<�O�k�wM�/��d����r�?�?�cx���P�CJ�p����-�gy�G��n�߱�j�_�nF4���Bϭ�ş]Ҁ�mD��D�r?���-�c����O�Q��S9��3{� DF~.�o	��5mhlm��3���G{�
�~���A|�y!Ѥ�7 q�������B}�N�I� f6j� �{e|�9��W��O�k����ѿ�N���8ke#��;��z�9����ܗ������>��5�������W����8f�ihƻ��p�Cؗ4'y�U-�ϟ��~����CO˩��Z��x�_���8��7~�J���.j,�Fgg�?�k6�DKG�ςOA�o��ܰ-�u`� �=E�� )�m��b��E�Qn���d�^}Y�I��T�/���ߋ���i�7۵���4�n����s�!�Zy�g�,qiE������9u.
�c����+pn��="ǜ��4@l�̮:���R��i�?�|�N���oc���"�*7���f��x43߯8:"-��XC}�x�hX�!��q)��̬�9�BaT��>\���v��O�o��!�����j�K��"��������A����n*94��
%��B�qq��]ґ΄WN�_��o�
С�O�'��W�����
$s.�h��R[Wc�h�����W����O�^\����o��У��4��U���gmD� lR����0��z2���4�y�D���ӗϢʴpYj���.��'�ڢ5Gl]*��կ}��&>��?���cV�X�o�P���%�)|q��X}�usFY#�"�Aḱ����G��C,҄~K�ݺ&�&Ӛ�����d��f3��� ���'*��$����b��ZL"�@��B�h
`�aQ��L��{zW�q4�Km=��v T�Ǐ��/^ډ.|�v��cq`P+R2��62}ux���j_��t^3��R�?BB�$�N����;i�f���P���|/[׎!�G j2�0���"}�q��L������*Nt�&ҩ4~��m�;�	��,�=%��)�i�x����$No�L%sO���oE�X��`7�֣	�ive�8X�}fVP8f<��P~�_�<3e�eY����&j�#B-i��Hv��� tV����H��y&<B��qH��U��B<�:wA���j�+Ŧ�}ų6�lh�HN��3x���qY��z"W�_?܍�>xڢOR8���v>����"#Zq0f�0��3Ԃ}�������_U�U�"
ł��щ����N2�����Ey��O�V����M���ܬ��>o �V�������Π˓֨yA��=(v�{�<B��[��.���cG1*t����E�����H~��E�$󝿂=�-��0��U���[x�ӈ�����眦�9�-���p��t�aDl@����I>/�������'�p�F���7I1���	�M�H$�P ^9v^\�=��h�j����*z�Ό�+0-(��� l��r|o�aQr��C��{�r�aL��߿���^.��k���+z�x�~��oA�CF�/��D�}��Q����䳼�n�6p���x$ #@Ԃp8��&�jj���yPh��a�L�������"������ˊ��S�LC�*��>G^F��b�1
�R����_���~����;���99�Y>�v&_�zB�o_$�����TsQ��������<�eE����1!n�Ψ��W"Z�	S4��HC�����ĿIU��.h_S�N0�HS�.������ ,���'�/�Q`mk2cmgRp�p��t���
�����f{睑Z��Ł��_����[�6cC��A���$���^��ʈ�E�	�tB�g�׳Gc��q���cssma�^�@<��C)�/�$�m��H��N���H�m�3��J�j���ȗ�a�Z ���j��@�4�C@�4�ڈz ~F\]G0T���j��ޣ��4�Ǿ�
~�Ϙ����1[m�%�4TUc|�<ڽ[�h6�{5J�Ϧ\\2�0���"��嵸�#�3۫�Z����Nd�\o��&�>3�8��Z^o)�="^�����4=���8�7��N6ͫ��1_�q��1qK��¢M����Y�RꩍD�`����h/"��Q�tv<M)���M�Ŗ�Ɔ��ԾP{��Ʊ�O�|N���9�J�ѧFƻ6ቾ�zX��WKlNϦ��d��x<�������P��p��T�X"�ʹ%ÃRO �_�vă�"�vb�4%ƛT��N� y}��8���<+G34���Ą�O��M $1	%��� j-����%�Mcο���M&m�E0��O]cj�_�mY�g�L�x2h̍��\-'����gpQ�;�w���+mg�8��b$q��#Z�0�v��t��p�qHNE��SSi��P��#��eR����f����&�	�C�lO�.�v
��Ez*��ڔ��9�AdV��#�+5�������XH���H��j��X�95�Z������x8��ED�Ƿ��˨�<�"����̓���}ݝ�P�R��9�)0v�ωƄD�>���)5��Ű766`ddt�����8JS��Jm
�:Gc���4Em����tF$=1�L�!t�y^jhT\h��;ڴ=�)����Y����x�Y�_�n����R1 ̪�3�4l�+jG_
x��GB�t��L�qa
��NA�J\B[�DR��;Ku�4������DF��
\X�l||L�.�P�|���3VzXK��Цp>�(�����=:~��FV�I����ȧ��@��,���.���U&�J��"�Nk�b�DS���-P>���ʏ����%�����"�0����QK�,�TJ(�ߡ�{�&�6��S���(.���IEV���ߥ�gE��.�O��-���|R�I{��d*��?ֺ�pF��+���ہۚίx"�2@��2Q�Ev>@�F26^�� S��d<a9�D��x<���_wvMMD�v�5w������t��d4J�����!���83b'�� @�Ietx>��Gp�J��_��A��+Z��h�Fl��[��ӖppnI�E[C�B[f�Ue���|�v�yq���+9	��:���(�P�C4ޤ	#m�&��'��kˑF;´�-��A��z���Dی�)`G���M4�c�X<~9�/x�cM�,{m����3����$��W��^�-�e�n�u��w:L� ���ؒ�/7�;�Kg����3dkZ��'�0�Û�u�1��tO�TC�� ��fΪl_��ŗ��Q){^�����w��IN� ��T�J�o;��Ǚ�JIl��Ԅ�h�^� b��#��ö�~�Ŀ�"�Z4 ��4'О���K&����7HP�v�.�NJ =p4ڥz��`0�B���*�������q�:�-'� �P8�C�s�h�}
�#���sF���x>��j�i��EЩ5�a���IAu����M텧87mq���!xjO��E�h/������d�f�Xݾ4�����(�(�[˘��Gj"��ǸD�� �*�?84�6��`N��zFl5KmS��g�X��������Bw	���DP[80P��3���$`��Б�w�抈z�h.�I[�O�֐؛��׵H5�@C�ܰ81���%0�CU-�R53��F״ TRCM�`�g���S�D@HS�I�6B]�B��%�sNEO�n5�OȨ�k�cs��⤦*e��A*#|����raH iI�+��|q�Sf-�zB�hɏ�����G�{R6j[j"��x���(omm����j)G���
�zE��`�S(HC�)��:�=v�.ٗ�zY�/��0R��%@)��` 5Ѯ0_VT:�M��dR4��X�X�9��)�`1��bG��,ְW�e٨�G1�
<0�[5q
�P�'����GC=#��6R��{���4R�IQs�m���x�B���E1��#o�����D�HCuu���pV��D+ŗ3��h�(6�V4ҭn[�b�<ґ���t˷���E¥U2�˂�T�BZ�jc5bi��
��ά-��F���¢0�����;��;IH˚L��3�1���I��S�z�i�j`<W-"�Q9'��6�Im!�Fuj��G(���P5��p�nK�"d��O r)�bf��u��h ��T������дPH9BAK85��1K�i�9yE��J�6�*�c�N4�� 0&r���&�E]Q�y��ΠN�����(5R�����ؘtd+8Ԝ�ۧݴ�a��h��)'ߊC�5�"]����n"+Q��:ڎP(�.-���נ���a���֠��[���I4Ɛ��[�O.�F�/5�#���hs��u~ã ��(�1�jAs���40u��ޮ��G0��qG{p��	�oʉ��֐�bW���kӴ,T(O���	�11�8� 1֠�HS�'Ϩ���l
����U.=-�*�}�ǥ�R�)q��9�&�ir�G�X;ʔ�ޱgM�Ҩ!�=� �~]}���˰0EX�l�WE���5*/o\�A���*yS���
�#��A*� ��]HP�ω- �G�^^yS������΄T�%Vj��*��Μ;�������5������z���3�nU��B@�!U.K��R@7�p��C�8� ��`��o��J#�����W�+�d�؝rҐ�����u�ܱ���qh�9^����l�a�.7��h�G�_���ҟ����@:_DsP\�=o��Yڍ�ZE���a
�F�Jga��L%�z������Ç��Qe:�l����Fc:�N"�C�u�X8.,][��U�)h�i��6�ǣ��Uv�՝YC�m��0��k�	�'Dg ]E$�� �97 ����
g+$��i6�]�L�Z_��S�c�x50tݻ3��t�}9!Hꢐ>gq�
�\�P�S�R��}�3�����L���mcj��\
�U���ziL�v�?'�x\z&˩y����
��R/o��P�|�!E��^�V��ț�Rx
��A� 7�L_�Z� �w5�t-M��-Z��(HeR�F�"P�δԤr�0:�uZ���4�R�w'}���wx~����QE�n�z=����c�:f�'z�sf('�]<U��������HPu�
x�*��.o��466��0�qn�n� �Q_Sp�H4��,���ѡ���5%/���2!�X�Ȝ�G�3M��؃`���9u'�'�c�c�	�,NsP���)�:�FqݡaC]=�y+�P�P�ʭ�(�+j���ΨE+�4<c}�7t�/�a��c��s��p�G�E~'�����r"�҈� �Vm�H/�@(�r6@ˊL�2�K�4���z<&��̪i���kinnq*7I���:UaD^/+���s5�Fv���D��NL���^����:?��}���d
@S%�N�if�	A�)����0Mg.�e<�AX
��*�Q�N��3#X�1��r���ys%����y8��h���<���ĘO���`v�ʙƜ䕮��,R��DQ8ܞo��v{?���kCɛg�[�^����6_JOP�|���r���SZ�J�)��<�����ߋh�cn҅-S �;NPiN�<��]]]z��\	�������<���a]g?�\J����Q�"�� � JN�P¦5���%�+��t'�I���D�~\��s�t�P�15��}N4^
�(���堤)�"��UҮ����v"Q�Q��U��j][R$��U�Z�*��k~|���9Q+�"�e�jGF��j�����x_$��r��e=5��Ԗ@i"�I�%������D�U\�ct��)�>�I��Xp��F�P��dՊ F�bԝNg'��1��Hy�-����eD��b�FJyoS�ے�Z�4_c08�5*L�8��B9����������Y�ö���mZtLz��(�&h�k�5��^P��r0�%����46�5��yw�V����;N�}lf�<E[NjA�ts�Amdފ{8G=0��b[�p��j�����[�� aCRhk\���]�7^b ���Y͈����髹�^�㺆��Й�-{J�jS�/-?-�iJ����f8��D�")Hg���15x,E���Q�p��9t1����p�12/�6��u/ȥ�%�D��Ϲ���?O�i�3�x]_�2٘V!0��bj��r��3��T2�Q(-9`N�!}�g�Z,gAOA��JQw҉��=�$:9�ZZZ��^�b)��<��xt�^�Y����y��c��l)������/s<�BT�{�<Ɲ��>���V�.+��̭s�Ӹ'�Ĵ���4x��<��0"��t<+zS�#RO�47ο���[�qn����ڦs�<��ץU������8�ꍹ%FTS�k�7%ߗ`�\��T
ȱ�ҭ�ɸ	-������1X��"W�(Ӎu\լ�.XN�X��u�qu���(|f��	Ig�*;9�2i�D�LR؜�rJN���	���7���r?�[����ʂ��Fp����L0Na`hL��`��X�/��[�w?�0+1�O�+�O2I��2e�����&�ޔfqa���pJ�l{2����$
I|�q�� 8�6�k�Ĕ�H��;2��ﶎ`m�3��'I��&��2����~���wQ�)�w)�Vf����s0���Q�Z���՚ �RЄ�Ù($}�δ��6�9'�ҍV@��_��,O�����Sg��&��|�c��un߉y�5��]W8�M�|+�ʍ1���َ)2rٕ�E] Fi>��򎨭x\G���X����Gl��bϣ��L��FJ"��zA��z��Q]�Y,:�}�9s�Ρ��y'�.M��}F�+VtiI#p��c��f�%E^���,n(F[�N���Ʃ;&f�m����VA�5���n GHo�t6x�Z�
�s�I�?�����h�	�U���	�v�T���::W,���9��N?+'�!644��uC�jze�gB��-�V%�q�ك��#��)2偄���yYF�h
�@��a�R�ؗr#h�p�Z�����5ï⏼a����|��W\�$j���rl�n=^,NV�w�g>%�NߧA�չ�)��hm�r����[�v�2{ �BvQ`�n�ӳ{U��ˇJ6��Ȩ����^�Iu�I��R]�3���f�<}M.�[�I�f�3�/C������TBsX��Е�B_\�d{]�3�Lô��8	I�G��. ��)�@kl ����>�ՅQ�9����~$ #Y��3�F�N�>����1O�삶�Ϲ�/abC�Lk3wcond�"3����p�
��e3�遷�E�D�1���3Xd�Tyj����1���؇�}Bc���8�E������g~�<�;P����ĬQ��И!��S�T���	G|�����̀���K7�\�
�&�Ĉ�Fk���y� �G#�t᠀�od�`R�T�Y�2�d:�Ύ���
}�Q6 ���94Es!3���Z5S�w	1]���5�vh?��	3��Oeq��1_�2
"�N(h�җv��[[e/�T�|�3u�s)�I��<�z����>�����1	Or1eG�r���[M�`XN��g�mK�{��f�"`d�'C�Zb�O�ސ.cXl����F�_�AW5���s̮(��j[�;�h#Ju#K���k��˧t
)[���Q���w��$�0Fs6^���9�o�e��C���W r��Z�%3*o�}����Ćj�n�&p*m��L��ⱏNZ�4G���?f8ف?/�y0�zr�,�U�:��S��L��as�M��%}�%��:7
�s��6�SƱ,����^��=��:t۽C�1��F�{a�rΖ��D��D�WTA�b-#T�Z����qnK���-st�<-��;�9�����
�j6�R{H찐V���)�	J���	�˥1�|Iъ��M�M�[V;k7>��b��k�,��e~!�9G�]̈��8f��_��{,�tJ�Y�=�;�¦DV�_��^�'zQ��b��Pޅ�Zέh�r�|�ђ=��g�t��E�5I2���-�5� �-��|=��|^6��l�hD��AU:�d�v<�i�D��	�eqC�T�j<�[�_����m���=�:�ݧ��rc��ʚ�bT�?9n������g �������n.���/v� /TFWlK��e��鎷����A$�w���'�)Q�ڒ�hL��q��=��8�wf�Y�i�=^7��1Y�6�s�<s�c�\�+�G�~�X����c-m���ͩ[y�������ţ(2cZ!(�w~`��\��*r���;�������u9S�\�I1ڟ2|ѫ�}`ŤeӖ���-��h0���MW¨i�ؘ��Ҟ�ŊC������ګ�*��6
���`:�6�R2��IN.π#��oҞ����6J�s�>�=��B�a��rn�fUp�^qu�����t}�Rے��'m�V��{�<��̿&w΍�wc\��h��j��̶vD|�Q/�h
�KS��C;�yu�; ���ᄌ���N�a���6���o��ճ(P�p2�w\3Ҳ$�Qn'��t6<bK��t��� b#�ȁFy>3�����`(�G�߭�!X|�_BK����ԋy��O��X� .k^�j�6���ـ᮪���^�������#q�V��V�*�-�q0�m��Ц��+�q2�Iy`���i݀�\��#w�.T�`���x!��R��f����і�|��(vG����+���ݺwO9�<�!�����i�
La�߬v����U���Ft��R֏?~H���wNܼ���&,<��#��YU����vҞ�hs�z=�x�|2H+9����G�9l�xe<-q�S'ŝ�9z�v����E����~<7���ni���!-��5�E�H}}N'�<�i�F�.l��κ�	q�v
UҖ\��G=-Rg<�o��Xy6��@U��>iG*�����[pϣ��{���-����C�±yykX�M��6��|}ϰ��ѳ����w�=+jqmgDwb[U�B�ϽЇ{{��ym���H3��+��i���gHm��yh�Z�ù�[+�3)��ڌ��7�{����N�3N�(�q���	4��\��Ӟ�w%�������.�6�'���C��m!}��]Sb�c��l��'4���o�"�1� ������#�R����9�:�V���)Z�6� ��?��w௶w����(O���D-v��SZ��l$p��I�,��^{n�ߌ��o`��Jj���XF)�B�L���>2��4W㌺ ��jA�!���:BhR����_ ���\A��#tH�O����Z #pg	�Q�AѪ����:<.�)��3��X�w}wԍ�/�}��ZO�ݘ�^�� s-an۵�j.W�wqVC��3w�x�d���1�0I����ʀڌOllR�a��&�����K�(��hA2���6���.�ݢ��[������-�q`���`���x;7�w���=���)s�����:�]\�$��4C�;�L��4�`c`�sjh?��Y>�N���w\�ӄ�쏩�#X�%
����e��#�m���R ���4�_�C�Kl�7,.6A���hk���2Ն@K4��C�O��}xמ{R�����='��.(��>����M��������(<�^1���8�/�:�*0W��(�J8`lBo��j	�&𐀒-!�Q�t�i�ig��U�v���L�\$:�v�ت�LA)lcį^��C0�Uf�d:�o����E ��`�_?0�^���E����q{��;��֥��ҍ��?���hط��5	�#�PP�b��7��g�������q�R�����g�lW��Β��������<��\����2�A����pk����}���H����m����K��H?�w�p� ��Uk�?Ule��=��Vq���V��G��p�-�p���%�b�?+�|��j�ls*�9&Z4�f�`ow�]��;n��ϼ-��`��q�y�߼���������t���`���-3E4�oG����[9���6�K����mm��]��}�V��X�l��)n�D�=q|"�g��6�g�
��E'9֘��2@��7���>�=|�}書.���ӧϗ�,�i�]7���Ŧ�����-���@��R��H?���kn������é��9���q�2�e��o�<���A��u�4��~�|^񼌊��4��>S���`h:��ʵ�$Sxl,���0t�j��jTNE�l��r+p#2�ۮ��o��WF瞟���!�]c��*���)���s�y�r���C&�ǁXO$$��ق���w���{^�`o1�����@@b���Aߖ��;�/㞽am�8���*�A��>���r�:���Jt��e��sֻ�%�`��+e�%wz�߁�E��۲AW�������ܸ�Tw
2�^{
�z9>�z_���y4����� :]q�zlԋOZ�15�`��9��f�KK��h}8g�/o�ۨFoh�[6�е�����V�.��< )7�'G�����"�/�P.�����1�wl ���ٸ>>����э�;��/�|}=
5�@m;�H+ܡ�n7���@ᔹ��m���M�&����&�$�m�o/�l�HK��m{ޡ���Rj�~#^�t}`K��.,��|���`P��@�1L��.	~Q�b��y�2��^b{�µ�L��7�]�ЛY̱�
�>W�tޣ-�Æ� V��	8�h��Q�3�F,�<�a��3/����O�o_W�_=���Am`��`�82�;v⡃Qб�oX����65񙷯T@ʭ?���Ѵj)� uE�h{q��z}�|�8���c�`
�������!�m���]�������p��<ߗP0��Ӄ���񻱹)��Oo�{�4��kk����s�~ܳ{tك��!<�_z�z���h�Ӄ���cjO��c���y�{�L���BU_�q�J\�:�o�#n�{/~���e�ª�KV��o�[�`�؟���e���n���l>����$n�Ϋ
���m��ɱ�&�x�;��1-Ƕ,!5�<�?W�-p���蝯�3P�F,�1wb�����ߟ�wH��G�n�_�1����H�/]~=۲$'�-�aM�3��;?:�t啑���h��*U�Ą�~0��D�x�2ް��ckK�l�¯mo��p�d�F�����g������ ;4������-���g4���wmY����o�pn��U$,��w��{����f��"N���s�iɲ��qՆzԉ�$��ʓ���*	 ����RxR�L������:V������t�Cg6+�}��>���ڌ�O�Q�-�jpٚ�'�t�	Ȝ�\���N��WGqH"oړ[���ٟ��?�X�8͆��E��e]�ӷ����8����)g�Npy���m���֖ 4��>���H9�SB5�vi'���p˿��7wh��^��rM�GE�Q4���b�����N$��ZN��XkY�y
1�wv����pzkWHtΈ{mC@m��=ޫn��u\^5����ژ�*7v��L�)`ɿ��YV��M�ޞ�Q����*�^����ӊ��}#i<{4>���fqo?*�����?�}̛2�OP���<�7��9�����ﾆ�jg�p"�v��ڇ?��C����a-�;Q�?��;/���S�r�A��\�,��Yf�,+@��I��)0���/\�F�7���ct���80��R[S�K��E�
(�Beqq�[r~YB^#6`4U�}	�4������p�xG����\zY��Sx._�,m�6<y$6io�om��>��R��Ŀ�R(���
�9n��iJ)���K�:�M�������W��(���`�yƔ���W:�+�$���LH��\o|2	Yv�q �,g~� tx�g�-��'/l��{L<��U|��61��j���AG�������8,6dH�.s-`����0.[QJ����e9i�� ����k����g4��ǽ���g���G%�G�����[��,c00�΋�](=Z5�+��g�\�}�x~��e��_v���S�7�������׮A<���=��L�Q�K5�3�9A��]H4cu���p66���k4z��v�-K@(L�߽� ���ͨzpǍ�🅺��7��t�C�� ��+_z�:�q@NpH0�s>dq�s�`�O�߃��F�g�q�i���~|��~˨M.�}��<I)���bV��M
���;�������
��xS�}��]k5%���[�4�BOi�ȁ�����p����,6���f����@q9�eAa��o��ߺ�]G=��wz���(p��3�RLP���kR1�y���4y�{��EF�ub�X_���<�Mח��3=1|_�GNh��F ���(L�Nd5���z����UT��j�i�c��<�rj�r�k�1�`{� Rn�R�M�b��0u	�K��ò�*���� )���Ms������& ˬ�	�2ko��ڛ�,�� @���ϑ��'�Z,m�J������,��9�	������c{��-4M=�X���q�Y�KZ����>��l�pN���=��T~�i��,���Y\`��	aņ����M�{CX��0�=���Z�7*'�������Tх�cFy���>��ˡ�	W�V]��5�jPtO> ��_�F��T?<����]'ԖY!�b|^.�
�6�����q>a����t:�zW
���ֆ�ǎ������LX������fz���������.>��o�r��=U*�{��TM#���a��^[��TN|,���r2=I|b��L}�ߙE�`�
�q�Pͼ����޲�U5u�8S1[�C����q�g��>�ti�<!}٦��4��=x�<���mYOF����:������ke���șA��!�]αG�����-���ݔ�6r.F�~h\�wi����;��'��S���O?��0��oHC�
&����+���z���)�5n��g�^��m�/��볻f�iƷ�f�x�J��kDS[�>�|��hjjDMMo�ō#���{�)RA���o"���(�qOd	g�0w܊�sC7�l��Ϩ����5rq�����������7�&��y|�|9V�����E�QWw�Z3�r�翅�3?
4��E;e�gӸQh���"�NՊ��i�����q��/���m�U{j���ѕ�{OoF[g|��O2����m]+�T?:2���g�J�Y�!�6��,,���1#1H�׉P�'�A�Uc�t'����	���
2������o��Fq����uHh_��Y��m�H�r��`���*:��{K��i<^߂�D�i9ݴ5��{F0QtOc�i��E����k:F����[׭�Em��5c�xa�	,�nG^n��?F����n+W����ܶ�y
�G�N�7��l^��uI_�d�T*�"��.}C���e�MT��t��jJߴ����P��7M�ς���v�Vw-
�)����+�}G���%� �n�gv���G�M����p��>`��m}r���|���U����"xc�	��Ow!�r����en��Vu��ʷnP՟����D,#�l �v���+NS>�'����G��-o|ƾ��ո����[@����vcx4��d^�}\e��vvW-��H�bry�pM~�=H>�| |���Z,5����V��>s|�|�#�#��#��N>Mm��&&�������	�O,ƾdd��'ta��x<���ʋw�ƠoU�m��j�����7ݨ�����|"ڋ����[8.B�N�dD���	EG@bI�EY긔s�Z4M�F�x������S��v�<׭�%�����r��m�Q��L/�<}���m�g����ӓ��"���.��D6gaz��㒾C#I�˨��JE��5���wd,�g�Oj��BNg��%�=��Q�.��7��d_��%L6�W��n�$ȩW�4s7��%�to���=��=��]�魘�Q��g�:[&Z�Ná2����y�0'�)}�S��,�,J@:}�B�x�oa��ޜ�R�D2+�Q�Ω}�\�,@��OM���K�Sw���O���,���Jk�~^�.��(��.�_����$r��͖/�ܛ&7�+��up2��~n���� NF��ګ����;�	��w���~t��xyna���2��ʵ^��l̈�)'�#�5�,aN?z(z\����ѻa��W����J�ɋm�_�u�Ǘ�غb���G�v�5��6ꓑ���]�.��_�#�������p�4��}EOз�jd7^����^���>ysf_n�ܷ�Jd6��������}�ҷ8Ó��H�o�ې�|w�?.��"��ן���_�Y��(��D�89/Ӹ����0�>mq��#�]_z������Bf�U8Ը^5`�����*؍�5eA�n������O��7(}��c�rފ#u+�ʥ���	H�҃��mͯ�Gj:�o���2`즵��Qn��/=ދs;ødU͢����FUƳ��������jϮY (��?ܫ���Y]�o4�W����r�B�5}1o_^;�E����� ����5�"��������Y���Ҹ����l)�ٶ!�� ّ����k/n>�YK8Y�<[��'��z���5oU�d[�C|�C�Y��>r�k���o�תkgkܫ���ŷ��T͉��$ ��F�2��&����\��FԳZ�=��ܞ;�bh�2uq��O���4��>vw�8��긜�����7�ó�u>!rN�K���XN$u���4:1�x���v�L+�����(u��Ws��4���W�񃗇���war����u���N|Bc�u�o6��K]�f6qy���<%����#y�����hL��$���F�y]/�{�E�j�o���Q��c�E^����_�ޑ:    IEND�B`�PK   ���X�B�>�  �'     jsons/user_defined.json�Z[o���+��NQ-����d+-�&vj7�C{cB�T()AN��ޡ$�r�OPѓD.���η3߬�M7_Wqz2ݮc�>Ĳ�c�Φ�c���n������������s{�=����MN�ho��	��v?4�W;}Y��������`�d�n�lZ�����(�{�<�ȕ�GX3eJa�����"�}[�6{��<���r˘D>z����R���:�"qŪ� �U����*�@�@�[��(r4����Y�.o���混���������e]6ӓo�z{��֫��z�,�MM�� �D�n]6_�[�D1������O[�T�2\m�
��Jt�u��~]-�
ôP�1#�����\�k��i�����.v\��M�φ�I�w�B3��/�r}���$>��>�&q��g=x��s-e6����V�_{V|�Z���p�mV��T���!��Y5u�7׷D!�cy1oö�����G�x]��� ܴ�r�=~��AYp�C$+!0�(��b�v�(�8��G�i�X��2�b�A!����S�:�z��uv?���=���QNM!�B����M��3���~{���E:��AM�0�Pxyq��o#b��,�˸��1Ld,+�u��QU�Hc�>���<�C�>��Ӡ�Jq�5\K��>(���$��c&���ÿO+��s�퓊�E���A���y�?�i�>�h^��E��'c���'A��^�Q�3a�4� �H���H��"4�YI�X���.ȑ��s��\�4�@���i�ҁ�%sa��HZ*֤Qr��D�i�>�v�v�J��9FI&�L��)�K9��]��-�����@�♨izс�%2Q��b�Kf�������D�)up�%�d��bB^�8�%rL;��]I-���[-�@R|���뽣PC�5�ͪ��]nw��Ĳ8���P�l�\�g H~x�i��j]�e�q����;wt�zRm�-��l[&�L��O0=,���뾸zS�?���*��w~���NC�`�!g� �5�;D�",0a3������h$1($n�B�F�\ĪLˈ�a)�K���f��qx��ӓrh�����CEnxņ�3\t���uHB��N�rq\D�+Gj�aW�Fa��r7(��#��/tǳ��$�0C=�i
f���=o�϶��F[���V�tBZ��v
�UrF��%�@�߳3ز�V���:l�g����t���u\N.#���7q=!x��G�y�|y�b!��u%2�Z$J�Q��v�KW�R���N�%ԫR#]Z
u���!k�#`D1�o��h[�0b�`[��b��w>��B
B������>����S�g�ZkÞ���P��f7��Xc�M@�3I����@����d:w�]h��G��.��h;,���<a�<ݙ�W��0�;�m��Cns�n���0��F�P�ʐ6�CR)�����'}q6y�l�vTF�1�Pye
�����"�5�e(=�g66�<2�)'>�����b�����T
>zY�2�P<��'�PD�z�x2:���A�U�
}̓���HœT.���b8�/$`*?'��]���ɪw�#!F���h9Ұ2�$�d�xEi�y}u��k��X��i8����(=i#�F�$�
䬳Rh�讏��V(��#����-��1��p�Ɍ<�H!��E��������5���i�(�vj���خ��d�V��ܕ^�:a˘�c�����_�_P?��/����Gdb=~/F�_���/N�-���+?��i:��_�s,��:�X�G��Cg��1q�`a�\�9k}�a��9�Hw.�G�3�8M�\K�3H}�c�$r���U[�6��Z��~&�w�z������3�18�d��U+�zrj7����V�
.R��X0d��H)J�)����+�[���
^"���K �@��¥�A��T$$��r�����kn�sX!OKce	u�quae�x�SEZ�=�� ���PUψ�`8퉁����{�ט>�p��S	�����dz���PK
   ���Xw�x5   r�                  cirkitFile.jsonPK
   ���X��(��8  �8  /             G   images/02932828-f6d4-4923-89fb-67d65ebd103a.pngPK
   ���XG�~��  � /             wY  images/0739a1b1-a163-452a-a325-ab452d55b136.pngPK
   ���XWC��)�  � /             N images/093f54e3-331f-4155-80d0-fca9fbcaa25c.pngPK
   ���XR�\"# � /             �� images/16f29068-8fa2-43fd-94bb-aa3b1aab738c.pngPK
   ���X�j�� 7q /             3 images/3afa6c98-60d7-4a37-9aec-be07fd386e0e.pngPK
   �x�X䏆ze� r& /             �� images/46a4a336-cec8-4b03-9de3-7f7682b07e1b.pngPK
   ���X����+  J  /             L� images/5644ca41-1cf6-484a-bb07-c2f9a6f5b19b.pngPK
   ���X��_8
  3
  /             � images/57489f55-55cc-4ea4-8258-f1cf3d9c722d.pngPK
   ���X	�\  \  /             I images/898ac7d1-13d0-4a1b-8b5c-ab7066f4327a.pngPK
   ���X�Ƚ׌  �  /             �. images/9185dcb2-65ea-4de0-8d42-42cedb1b5634.pngPK
   ���X$7h�!  �!  /             �7 images/c6364832-c854-438f-b38b-75bf2a0cd33f.pngPK
   ���X~��a� ٮ /             Z images/dc707dc6-8489-41bb-a5bc-77a0670f90d6.pngPK
   ���XP��/�  ǽ  /             � images/f42d805d-3c79-4d19-85d7-77e6ec425ca7.pngPK
   �x�XQ//�@  �?  /             � images/f7eed1a5-74ac-45f9-b2e1-80b6b3a4cd0f.pngPK
   ���X�B�>�  �'               ^ jsons/user_defined.jsonPK      �  �	   